<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.80168">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Campo Mourão" name="Torneio Regional da 2ª Região (Pré-Mirim/Sênior)" course="SCM" deadline="2025-04-21" entrystartdate="2025-04-14" entrytype="INVITATION" hostclub="Fundação de Esportes de Campo Mourão" hostclub.url="https://campomourao.atende.net/subportal/fundacao-de-esportes" number="39785" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/newInterface/eventos/39785/" startmethod="1" timing="AUTOMATIC" touchpad="ONESIDE" masters="F" withdrawuntil="2025-04-24" state="PR" nation="BRA" hytek.courseorder="S">
      <AGEDATE value="2025-01-01" type="YEAR" />
      <POOL name="Estádio Municipal Roberto Brzezinski" lanemin="1" lanemax="6" />
      <FACILITY city="Campo Mourão" name="Estádio Municipal Roberto Brzezinski" nation="BRA" state="PR" street="Av. Comendador Norberto Marcondes, 286" street2="Centro" zip="87302-060" />
      <POINTTABLE pointtableid="3017" name="AQUA Point Scoring" version="2024" />
      <FEES>
        <FEE currency="BRL" type="LATEENTRY.INDIVIDUAL" value="2800" />
        <FEE currency="BRL" type="LATEENTRY.RELAY" value="11200" />
      </FEES>
      <QUALIFY from="2024-04-26" until="2025-04-25" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99252-0598" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99252-0598" street="Avenida do Batel, 1230" street2="Sala 202" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2025-04-26" daytime="09:15" endtime="12:43" number="1" officialmeeting="08:30" teamleadermeeting="09:00" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="1060" daytime="09:16" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1061" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11619" />
                    <RANKING order="2" place="2" resultid="11506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11277" />
                    <RANKING order="2" place="2" resultid="11695" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1063" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10846" />
                    <RANKING order="2" place="2" resultid="10852" />
                    <RANKING order="3" place="3" resultid="10943" />
                    <RANKING order="4" place="4" resultid="11417" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1064" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1065" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10912" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1067" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11722" daytime="09:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11723" daytime="09:20" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1068" daytime="09:24" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1069" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11267" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11247" />
                    <RANKING order="2" place="2" resultid="11428" />
                    <RANKING order="3" place="3" resultid="11340" />
                    <RANKING order="4" place="4" resultid="11129" />
                    <RANKING order="5" place="5" resultid="11690" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10873" />
                    <RANKING order="2" place="2" resultid="11306" />
                    <RANKING order="3" place="3" resultid="11360" />
                    <RANKING order="4" place="4" resultid="11262" />
                    <RANKING order="5" place="5" resultid="11635" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10867" />
                    <RANKING order="2" place="2" resultid="11412" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1073" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11311" />
                    <RANKING order="2" place="2" resultid="11442" />
                    <RANKING order="3" place="3" resultid="10926" />
                    <RANKING order="4" place="-1" resultid="11239" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1074" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="11235" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1075" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11724" daytime="09:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11725" daytime="09:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11726" daytime="09:30" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1076" daytime="09:34" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1077" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="1078" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11035" />
                    <RANKING order="2" place="2" resultid="11212" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1079" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1080" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11479" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11727" daytime="09:34" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1081" daytime="09:38" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1082" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11085" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1083" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11060" />
                    <RANKING order="2" place="2" resultid="11483" />
                    <RANKING order="3" place="3" resultid="11119" />
                    <RANKING order="4" place="4" resultid="11012" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1084" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11291" />
                    <RANKING order="2" place="2" resultid="11350" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1085" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11031" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11728" daytime="09:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11729" daytime="09:44" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1086" daytime="09:48" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1087" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11394" />
                    <RANKING order="2" place="2" resultid="10989" />
                    <RANKING order="3" place="3" resultid="11331" />
                    <RANKING order="4" place="4" resultid="11448" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1088" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11296" />
                    <RANKING order="2" place="2" resultid="11705" />
                    <RANKING order="3" place="3" resultid="11711" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1089" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11301" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1090" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1091" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1092" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1093" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11730" daytime="09:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11731" daytime="09:52" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1094" daytime="09:58" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1095" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11423" />
                    <RANKING order="2" place="2" resultid="11345" />
                    <RANKING order="3" place="3" resultid="10891" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1096" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10888" />
                    <RANKING order="2" place="2" resultid="11286" />
                    <RANKING order="3" place="3" resultid="11272" />
                    <RANKING order="4" place="4" resultid="10856" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1097" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11389" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10881" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1099" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11240" />
                    <RANKING order="2" place="-1" resultid="10884" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1100" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10842" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1101" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11732" daytime="09:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11733" daytime="10:02" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1102" daytime="10:06" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1103" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11552" />
                    <RANKING order="2" place="2" resultid="11543" />
                    <RANKING order="3" place="-1" resultid="11532" />
                    <RANKING order="4" place="-1" resultid="11535" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1104" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11502" />
                    <RANKING order="2" place="2" resultid="11096" />
                    <RANKING order="3" place="3" resultid="11560" />
                    <RANKING order="4" place="4" resultid="11198" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1105" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11474" />
                    <RANKING order="2" place="2" resultid="11373" />
                    <RANKING order="3" place="3" resultid="10862" />
                    <RANKING order="4" place="4" resultid="11624" />
                    <RANKING order="5" place="-1" resultid="11520" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1106" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11489" />
                    <RANKING order="2" place="2" resultid="10993" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11734" daytime="10:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11735" daytime="10:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11736" daytime="10:12" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1107" daytime="10:14" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1108" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11086" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1109" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11355" />
                    <RANKING order="2" place="2" resultid="11061" />
                    <RANKING order="3" place="3" resultid="11013" />
                    <RANKING order="4" place="4" resultid="11556" />
                    <RANKING order="5" place="5" resultid="11041" />
                    <RANKING order="6" place="6" resultid="11539" />
                    <RANKING order="7" place="7" resultid="11188" />
                    <RANKING order="8" place="8" resultid="11549" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1110" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11115" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1111" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11320" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11737" daytime="10:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11738" daytime="10:16" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1112" daytime="10:18" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1113" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11081" />
                    <RANKING order="2" place="2" resultid="11325" />
                    <RANKING order="3" place="3" resultid="10997" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1114" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11255" />
                    <RANKING order="2" place="2" resultid="11377" />
                    <RANKING order="3" place="3" resultid="11464" />
                    <RANKING order="4" place="4" resultid="10957" />
                    <RANKING order="5" place="5" resultid="10969" />
                    <RANKING order="6" place="6" resultid="10992" />
                    <RANKING order="7" place="-1" resultid="11469" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1115" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10965" />
                    <RANKING order="2" place="2" resultid="11618" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1116" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10949" />
                    <RANKING order="2" place="2" resultid="11335" />
                    <RANKING order="3" place="3" resultid="11710" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1117" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11700" />
                    <RANKING order="2" place="2" resultid="10940" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1118" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1119" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11228" />
                    <RANKING order="2" place="2" resultid="11133" />
                    <RANKING order="3" place="3" resultid="10922" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1120" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1121" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11589" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11739" daytime="10:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11740" daytime="10:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11741" daytime="10:26" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11742" daytime="10:28" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1122" daytime="10:32" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1123" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11050" />
                    <RANKING order="2" place="2" resultid="11349" />
                    <RANKING order="3" place="3" resultid="11008" />
                    <RANKING order="4" place="4" resultid="11367" />
                    <RANKING order="5" place="5" resultid="11566" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1124" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11280" />
                    <RANKING order="2" place="-1" resultid="10978" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1125" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10982" />
                    <RANKING order="2" place="2" resultid="11404" />
                    <RANKING order="3" place="3" resultid="11627" />
                    <RANKING order="4" place="4" resultid="10986" />
                    <RANKING order="5" place="5" resultid="11266" />
                    <RANKING order="6" place="6" resultid="11453" />
                    <RANKING order="7" place="7" resultid="11576" />
                    <RANKING order="8" place="8" resultid="11648" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11436" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1127" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1128" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1129" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10915" />
                    <RANKING order="2" place="2" resultid="10877" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1130" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11605" />
                    <RANKING order="2" place="2" resultid="11103" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1131" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10953" />
                    <RANKING order="2" place="2" resultid="11581" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11743" daytime="10:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11744" daytime="10:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11745" daytime="10:38" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11746" daytime="10:42" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11874" daytime="10:44" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1132" daytime="11:04" gender="F" number="11" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1133" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11192" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1134" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11036" />
                    <RANKING order="2" place="2" resultid="11065" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1135" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11458" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1136" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11510" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11747" daytime="11:04" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1137" daytime="11:06" gender="M" number="12" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1138" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11125" />
                    <RANKING order="2" place="2" resultid="11528" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1139" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11120" />
                    <RANKING order="2" place="2" resultid="11091" />
                    <RANKING order="3" place="-1" resultid="11498" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1140" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1141" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11321" />
                    <RANKING order="2" place="2" resultid="11021" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11748" daytime="11:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11749" daytime="11:08" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1142" daytime="11:12" gender="F" number="13" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1143" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11075" />
                    <RANKING order="2" place="-1" resultid="11080" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1144" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11045" />
                    <RANKING order="2" place="2" resultid="11478" />
                    <RANKING order="3" place="3" resultid="11463" />
                    <RANKING order="4" place="-1" resultid="11468" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1145" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11407" />
                    <RANKING order="2" place="2" resultid="11330" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1146" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11276" />
                    <RANKING order="2" place="2" resultid="11295" />
                    <RANKING order="3" place="3" resultid="11493" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1147" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10851" />
                    <RANKING order="2" place="2" resultid="11300" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1148" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10908" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1149" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10911" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1151" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11750" daytime="11:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11751" daytime="11:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11752" daytime="11:16" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1152" daytime="11:20" gender="M" number="14" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1153" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11002" />
                    <RANKING order="2" place="2" resultid="11290" />
                    <RANKING order="3" place="3" resultid="11070" />
                    <RANKING order="4" place="4" resultid="11007" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1154" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11030" />
                    <RANKING order="2" place="-1" resultid="11025" />
                    <RANKING order="3" place="-1" resultid="11055" />
                    <RANKING order="4" place="-1" resultid="10977" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1155" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11315" />
                    <RANKING order="2" place="2" resultid="11403" />
                    <RANKING order="3" place="3" resultid="11422" />
                    <RANKING order="4" place="4" resultid="11344" />
                    <RANKING order="5" place="-1" resultid="11571" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1156" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11427" />
                    <RANKING order="2" place="2" resultid="11271" />
                    <RANKING order="3" place="3" resultid="11432" />
                    <RANKING order="4" place="4" resultid="11339" />
                    <RANKING order="5" place="5" resultid="11285" />
                    <RANKING order="6" place="6" resultid="11640" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1157" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10872" />
                    <RANKING order="2" place="2" resultid="11251" />
                    <RANKING order="3" place="3" resultid="11261" />
                    <RANKING order="4" place="4" resultid="11359" />
                    <RANKING order="5" place="5" resultid="11305" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1158" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10919" />
                    <RANKING order="2" place="2" resultid="11596" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1159" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11310" />
                    <RANKING order="2" place="2" resultid="10936" />
                    <RANKING order="3" place="3" resultid="11441" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1160" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10841" />
                    <RANKING order="2" place="2" resultid="10902" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1161" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11232" />
                    <RANKING order="2" place="2" resultid="11600" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11753" daytime="11:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11754" daytime="11:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11755" daytime="11:26" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11756" daytime="11:28" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11757" daytime="11:30" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11758" daytime="11:32" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1162" daytime="11:36" gender="F" number="15" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1163" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11395" />
                    <RANKING order="2" place="2" resultid="11408" />
                    <RANKING order="3" place="3" resultid="11449" />
                    <RANKING order="4" place="4" resultid="11620" />
                    <RANKING order="5" place="5" resultid="11507" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1164" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11706" />
                    <RANKING order="2" place="2" resultid="10946" />
                    <RANKING order="3" place="3" resultid="11494" />
                    <RANKING order="4" place="4" resultid="10950" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1165" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11701" />
                    <RANKING order="2" place="2" resultid="11632" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1166" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1167" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10905" />
                    <RANKING order="2" place="2" resultid="10923" />
                    <RANKING order="3" place="3" resultid="11134" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1168" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="11111" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1169" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11590" />
                    <RANKING order="2" place="2" resultid="11683" />
                    <RANKING order="3" place="3" resultid="11100" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11759" daytime="11:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11760" daytime="11:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11761" daytime="11:38" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1170" daytime="11:40" gender="M" number="16" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1171" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10974" />
                    <RANKING order="2" place="2" resultid="11454" />
                    <RANKING order="3" place="3" resultid="11628" />
                    <RANKING order="4" place="4" resultid="10962" />
                    <RANKING order="5" place="5" resultid="11017" />
                    <RANKING order="6" place="6" resultid="10892" />
                    <RANKING order="7" place="7" resultid="11649" />
                    <RANKING order="8" place="8" resultid="11644" />
                    <RANKING order="9" place="9" resultid="11577" />
                    <RANKING order="10" place="10" resultid="11572" />
                    <RANKING order="11" place="-1" resultid="11653" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1172" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11437" />
                    <RANKING order="2" place="2" resultid="11130" />
                    <RANKING order="3" place="3" resultid="10857" />
                    <RANKING order="4" place="4" resultid="11691" />
                    <RANKING order="5" place="5" resultid="11399" />
                    <RANKING order="6" place="6" resultid="11641" />
                    <RANKING order="7" place="7" resultid="11592" />
                    <RANKING order="8" place="8" resultid="11515" />
                    <RANKING order="9" place="-1" resultid="10933" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1173" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11244" />
                    <RANKING order="2" place="2" resultid="10930" />
                    <RANKING order="3" place="3" resultid="11636" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1174" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10868" />
                    <RANKING order="2" place="2" resultid="11609" />
                    <RANKING order="3" place="3" resultid="11597" />
                    <RANKING order="4" place="4" resultid="11661" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1175" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11107" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1176" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11606" />
                    <RANKING order="2" place="-1" resultid="11104" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1177" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11601" />
                    <RANKING order="2" place="2" resultid="11680" />
                    <RANKING order="3" place="3" resultid="11582" />
                    <RANKING order="4" place="4" resultid="11614" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11762" daytime="11:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11763" daytime="11:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11764" daytime="11:44" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11765" daytime="11:46" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11766" daytime="11:48" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11767" daytime="11:48" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1178" daytime="11:50" gender="F" number="17" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1179" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11551" />
                    <RANKING order="2" place="2" resultid="11193" />
                    <RANKING order="3" place="3" resultid="11542" />
                    <RANKING order="4" place="-1" resultid="11531" />
                    <RANKING order="5" place="-1" resultid="11534" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1180" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11213" />
                    <RANKING order="2" place="2" resultid="11559" />
                    <RANKING order="3" place="3" resultid="11197" />
                    <RANKING order="4" place="4" resultid="11672" />
                    <RANKING order="5" place="5" resultid="11066" />
                    <RANKING order="6" place="6" resultid="11095" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1181" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11459" />
                    <RANKING order="2" place="2" resultid="11326" />
                    <RANKING order="3" place="3" resultid="11473" />
                    <RANKING order="4" place="4" resultid="10998" />
                    <RANKING order="5" place="5" resultid="11076" />
                    <RANKING order="6" place="6" resultid="11519" />
                    <RANKING order="7" place="7" resultid="10861" />
                    <RANKING order="8" place="8" resultid="11372" />
                    <RANKING order="9" place="9" resultid="11657" />
                    <RANKING order="10" place="10" resultid="11623" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1182" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11511" />
                    <RANKING order="2" place="2" resultid="11046" />
                    <RANKING order="3" place="3" resultid="11256" />
                    <RANKING order="4" place="4" resultid="11378" />
                    <RANKING order="5" place="5" resultid="10958" />
                    <RANKING order="6" place="6" resultid="11488" />
                    <RANKING order="7" place="7" resultid="10970" />
                    <RANKING order="8" place="8" resultid="11676" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11768" daytime="11:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11769" daytime="11:54" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11770" daytime="11:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11771" daytime="11:56" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11772" daytime="11:58" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1183" daytime="12:00" gender="M" number="18" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1184" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11124" />
                    <RANKING order="2" place="2" resultid="11527" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1185" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11354" />
                    <RANKING order="2" place="2" resultid="11484" />
                    <RANKING order="3" place="3" resultid="11040" />
                    <RANKING order="4" place="4" resultid="11090" />
                    <RANKING order="5" place="5" resultid="11538" />
                    <RANKING order="6" place="6" resultid="11555" />
                    <RANKING order="7" place="7" resultid="11187" />
                    <RANKING order="8" place="8" resultid="11548" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11003" />
                    <RANKING order="2" place="2" resultid="11051" />
                    <RANKING order="3" place="3" resultid="11071" />
                    <RANKING order="4" place="4" resultid="11567" />
                    <RANKING order="5" place="5" resultid="11368" />
                    <RANKING order="6" place="-1" resultid="11114" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1187" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11281" />
                    <RANKING order="2" place="2" resultid="11020" />
                    <RANKING order="3" place="3" resultid="11026" />
                    <RANKING order="4" place="4" resultid="11668" />
                    <RANKING order="5" place="5" resultid="11056" />
                    <RANKING order="6" place="6" resultid="11664" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11773" daytime="12:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11774" daytime="12:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11775" daytime="12:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11776" daytime="12:06" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1188" daytime="12:08" gender="F" number="19" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1189" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1190" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11696" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1191" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10847" />
                    <RANKING order="2" place="2" resultid="11418" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1192" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1193" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1194" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1195" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11777" daytime="12:08" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1196" daytime="12:20" gender="M" number="20" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1197" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11316" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1198" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1199" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11390" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1200" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11413" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1201" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1202" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1203" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11585" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11778" daytime="12:20" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="11880" daytime="12:32" gender="F" number="98" order="22" round="TIMETRIAL" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11881" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="11882" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="11883" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="11884" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="11885" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11897" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11886" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="11887" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11896" daytime="12:32" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="11888" daytime="12:38" gender="M" number="99" order="23" round="TIMETRIAL" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11889" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="11890" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11899" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="11891" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="11892" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="11893" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="11894" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="11895" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11898" daytime="12:38" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2025-04-26" daytime="15:45" endtime="19:59" number="2" officialmeeting="15:00" teamleadermeeting="15:30" warmupfrom="14:30" warmupuntil="15:30">
          <EVENTS>
            <EVENT eventid="1204" daytime="15:46" gender="F" number="21" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1205" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11077" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1206" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11471" />
                    <RANKING order="2" place="2" resultid="11481" />
                    <RANKING order="3" place="3" resultid="11466" />
                    <RANKING order="4" place="4" resultid="10995" />
                    <RANKING order="5" place="5" resultid="10972" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1207" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11410" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1208" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11698" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1209" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10849" />
                    <RANKING order="2" place="2" resultid="11303" />
                    <RANKING order="3" place="3" resultid="11420" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1210" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1211" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1212" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1213" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11779" daytime="15:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11780" daytime="15:52" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1214" daytime="16:00" gender="M" number="22" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1215" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11293" />
                    <RANKING order="2" place="2" resultid="11352" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1216" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11023" />
                    <RANKING order="2" place="2" resultid="11058" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1217" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11318" />
                    <RANKING order="2" place="2" resultid="10984" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1218" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11342" />
                    <RANKING order="2" place="2" resultid="11430" />
                    <RANKING order="3" place="3" resultid="11693" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1219" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11308" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1220" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11415" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1221" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11313" />
                    <RANKING order="2" place="2" resultid="10879" />
                    <RANKING order="3" place="3" resultid="10938" />
                    <RANKING order="4" place="4" resultid="10928" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1222" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1223" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11587" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11781" daytime="16:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11782" daytime="16:08" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11783" daytime="16:14" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1224" daytime="16:22" gender="F" number="23" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1225" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11174" />
                    <RANKING order="2" place="2" resultid="11184" />
                    <RANKING order="3" place="3" resultid="11164" />
                    <RANKING order="4" place="4" resultid="11154" />
                    <RANKING order="5" place="5" resultid="11159" />
                    <RANKING order="6" place="6" resultid="11209" />
                    <RANKING order="7" place="7" resultid="11149" />
                    <RANKING order="8" place="8" resultid="11546" />
                    <RANKING order="9" place="9" resultid="11204" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11784" daytime="16:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11785" daytime="16:24" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1226" daytime="16:26" gender="M" number="24" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1227" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11143" />
                    <RANKING order="2" place="2" resultid="11223" />
                    <RANKING order="3" place="3" resultid="11178" />
                    <RANKING order="4" place="4" resultid="11564" />
                    <RANKING order="5" place="5" resultid="11138" />
                    <RANKING order="6" place="6" resultid="11218" />
                    <RANKING order="7" place="7" resultid="11168" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11786" daytime="16:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11787" daytime="16:28" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1228" daytime="16:30" gender="F" number="25" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1229" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11327" />
                    <RANKING order="2" place="2" resultid="11461" />
                    <RANKING order="3" place="3" resultid="11374" />
                    <RANKING order="4" place="4" resultid="11475" />
                    <RANKING order="5" place="5" resultid="10864" />
                    <RANKING order="6" place="6" resultid="11522" />
                    <RANKING order="7" place="-1" resultid="10999" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1230" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11048" />
                    <RANKING order="2" place="2" resultid="11513" />
                    <RANKING order="3" place="3" resultid="11258" />
                    <RANKING order="4" place="4" resultid="11491" />
                    <RANKING order="5" place="-1" resultid="10971" />
                    <RANKING order="6" place="-1" resultid="10959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1231" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11397" />
                    <RANKING order="2" place="2" resultid="11451" />
                    <RANKING order="3" place="3" resultid="10990" />
                    <RANKING order="4" place="4" resultid="11332" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1232" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11708" />
                    <RANKING order="2" place="2" resultid="11297" />
                    <RANKING order="3" place="3" resultid="11712" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1233" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11302" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1234" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1235" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10906" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1236" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1237" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11788" daytime="16:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11789" daytime="16:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11790" daytime="16:36" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11791" daytime="16:38" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1238" daytime="16:42" gender="M" number="26" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1239" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11004" />
                    <RANKING order="2" place="2" resultid="11116" />
                    <RANKING order="3" place="3" resultid="11010" />
                    <RANKING order="4" place="4" resultid="11369" />
                    <RANKING order="5" place="5" resultid="11525" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1240" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11022" />
                    <RANKING order="2" place="2" resultid="11028" />
                    <RANKING order="3" place="3" resultid="11057" />
                    <RANKING order="4" place="4" resultid="11033" />
                    <RANKING order="5" place="-1" resultid="11322" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1241" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10963" />
                    <RANKING order="2" place="2" resultid="11424" />
                    <RANKING order="3" place="3" resultid="11346" />
                    <RANKING order="4" place="4" resultid="10894" />
                    <RANKING order="5" place="5" resultid="11646" />
                    <RANKING order="6" place="6" resultid="11655" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1242" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11273" />
                    <RANKING order="2" place="2" resultid="10934" />
                    <RANKING order="3" place="3" resultid="10889" />
                    <RANKING order="4" place="4" resultid="11287" />
                    <RANKING order="5" place="5" resultid="11401" />
                    <RANKING order="6" place="6" resultid="11517" />
                    <RANKING order="7" place="-1" resultid="10859" />
                    <RANKING order="8" place="-1" resultid="11594" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1243" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11391" />
                    <RANKING order="2" place="2" resultid="11638" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1244" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10882" />
                    <RANKING order="2" place="2" resultid="11611" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1245" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11241" />
                    <RANKING order="2" place="2" resultid="11109" />
                    <RANKING order="3" place="3" resultid="10927" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1246" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10843" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1247" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11616" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11792" daytime="16:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11793" daytime="16:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11794" daytime="16:48" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11795" daytime="16:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11796" daytime="16:54" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11797" daytime="16:56" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1248" daytime="16:58" gender="F" number="27" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1249" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11195" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1250" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11215" />
                    <RANKING order="2" place="2" resultid="11200" />
                    <RANKING order="3" place="3" resultid="11674" />
                    <RANKING order="4" place="4" resultid="11068" />
                    <RANKING order="5" place="5" resultid="11098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1251" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11083" />
                    <RANKING order="2" place="2" resultid="11476" />
                    <RANKING order="3" place="3" resultid="11078" />
                    <RANKING order="4" place="4" resultid="11625" />
                    <RANKING order="5" place="5" resultid="11659" />
                    <RANKING order="6" place="-1" resultid="11375" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1252" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11380" />
                    <RANKING order="2" place="-1" resultid="11678" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11798" daytime="16:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11799" daytime="17:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11800" daytime="17:04" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1253" daytime="17:06" gender="M" number="28" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1254" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11127" />
                    <RANKING order="2" place="2" resultid="11529" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1255" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11365" />
                    <RANKING order="2" place="2" resultid="11486" />
                    <RANKING order="3" place="3" resultid="11043" />
                    <RANKING order="4" place="4" resultid="11093" />
                    <RANKING order="5" place="5" resultid="11190" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1256" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11569" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1257" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11283" />
                    <RANKING order="2" place="2" resultid="11670" />
                    <RANKING order="3" place="3" resultid="11666" />
                    <RANKING order="4" place="-1" resultid="10980" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11801" daytime="17:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11802" daytime="17:10" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1258" daytime="17:12" gender="F" number="29" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11714" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11158" />
                    <RANKING order="2" place="2" resultid="11163" />
                    <RANKING order="3" place="3" resultid="11183" />
                    <RANKING order="4" place="4" resultid="11173" />
                    <RANKING order="5" place="5" resultid="11153" />
                    <RANKING order="6" place="6" resultid="11148" />
                    <RANKING order="7" place="7" resultid="11208" />
                    <RANKING order="8" place="8" resultid="11203" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11803" daytime="17:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11804" daytime="17:14" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1260" daytime="17:16" gender="M" number="30" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11715" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11179" />
                    <RANKING order="2" place="2" resultid="11687" />
                    <RANKING order="3" place="3" resultid="11139" />
                    <RANKING order="4" place="4" resultid="11169" />
                    <RANKING order="5" place="5" resultid="11219" />
                    <RANKING order="6" place="6" resultid="11144" />
                    <RANKING order="7" place="7" resultid="11224" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11805" daytime="17:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11806" daytime="17:18" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1262" daytime="17:20" gender="F" number="31" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1263" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10967" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1264" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11336" />
                    <RANKING order="2" place="2" resultid="11713" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1265" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10854" />
                    <RANKING order="2" place="2" resultid="11703" />
                    <RANKING order="3" place="3" resultid="10941" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1266" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1267" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11229" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1268" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1269" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11807" daytime="17:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11808" daytime="17:26" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1270" daytime="17:30" gender="M" number="32" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1271" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11405" />
                    <RANKING order="2" place="2" resultid="11268" />
                    <RANKING order="3" place="3" resultid="11579" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1272" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11439" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1273" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1274" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1275" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10916" />
                    <RANKING order="2" place="2" resultid="10885" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1276" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11607" />
                    <RANKING order="2" place="-1" resultid="11236" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1277" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10955" />
                    <RANKING order="2" place="2" resultid="11681" />
                    <RANKING order="3" place="3" resultid="11583" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11809" daytime="17:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11810" daytime="17:34" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1278" daytime="17:38" gender="F" number="33" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1279" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="11409" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1280" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11278" />
                    <RANKING order="2" place="2" resultid="11298" />
                    <RANKING order="3" place="3" resultid="11697" />
                    <RANKING order="4" place="-1" resultid="11446" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1281" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1282" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1283" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1284" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1285" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11812" daytime="17:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11871" daytime="17:44" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1286" daytime="17:48" gender="M" number="34" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1287" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11425" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1288" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11249" />
                    <RANKING order="2" place="2" resultid="11274" />
                    <RANKING order="3" place="3" resultid="11433" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1289" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10875" />
                    <RANKING order="2" place="2" resultid="11252" />
                    <RANKING order="3" place="3" resultid="11263" />
                    <RANKING order="4" place="4" resultid="11361" />
                    <RANKING order="5" place="-1" resultid="11392" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1290" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10870" />
                    <RANKING order="2" place="2" resultid="10920" />
                    <RANKING order="3" place="3" resultid="11414" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1291" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11312" />
                    <RANKING order="2" place="2" resultid="11444" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1292" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10844" />
                    <RANKING order="2" place="2" resultid="10903" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1293" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11586" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11813" daytime="17:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11814" daytime="17:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11815" daytime="17:56" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1294" daytime="18:00" gender="F" number="35" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11716" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11160" />
                    <RANKING order="2" place="2" resultid="11185" />
                    <RANKING order="3" place="3" resultid="11165" />
                    <RANKING order="4" place="4" resultid="11175" />
                    <RANKING order="5" place="5" resultid="11150" />
                    <RANKING order="6" place="6" resultid="11155" />
                    <RANKING order="7" place="7" resultid="11210" />
                    <RANKING order="8" place="8" resultid="11205" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11816" daytime="18:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11817" daytime="18:02" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1296" daytime="18:04" gender="M" number="36" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11717" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11180" />
                    <RANKING order="2" place="2" resultid="11140" />
                    <RANKING order="3" place="3" resultid="11145" />
                    <RANKING order="4" place="4" resultid="11225" />
                    <RANKING order="5" place="5" resultid="11220" />
                    <RANKING order="6" place="6" resultid="11170" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11818" daytime="18:04" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1298" daytime="18:06" gender="F" number="37" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1299" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11194" />
                    <RANKING order="2" place="-1" resultid="11536" />
                    <RANKING order="3" place="-1" resultid="11553" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1300" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11038" />
                    <RANKING order="2" place="2" resultid="11214" />
                    <RANKING order="3" place="3" resultid="11561" />
                    <RANKING order="4" place="4" resultid="11504" />
                    <RANKING order="5" place="5" resultid="11199" />
                    <RANKING order="6" place="6" resultid="11673" />
                    <RANKING order="7" place="7" resultid="11067" />
                    <RANKING order="8" place="8" resultid="11097" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1301" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11460" />
                    <RANKING order="2" place="2" resultid="10863" />
                    <RANKING order="3" place="3" resultid="11521" />
                    <RANKING order="4" place="4" resultid="11658" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1302" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11047" />
                    <RANKING order="2" place="2" resultid="11512" />
                    <RANKING order="3" place="3" resultid="11257" />
                    <RANKING order="4" place="4" resultid="11480" />
                    <RANKING order="5" place="5" resultid="11470" />
                    <RANKING order="6" place="6" resultid="11465" />
                    <RANKING order="7" place="7" resultid="10994" />
                    <RANKING order="8" place="8" resultid="11677" />
                    <RANKING order="9" place="-1" resultid="11490" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11819" daytime="18:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11820" daytime="18:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11821" daytime="18:12" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11822" daytime="18:16" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1303" daytime="18:18" gender="M" number="38" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1304" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11088" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1305" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11357" />
                    <RANKING order="2" place="2" resultid="11063" />
                    <RANKING order="3" place="3" resultid="11122" />
                    <RANKING order="4" place="4" resultid="11042" />
                    <RANKING order="5" place="5" resultid="11015" />
                    <RANKING order="6" place="6" resultid="11540" />
                    <RANKING order="7" place="7" resultid="11189" />
                    <RANKING order="8" place="-1" resultid="11500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1306" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11052" />
                    <RANKING order="2" place="2" resultid="11072" />
                    <RANKING order="3" place="3" resultid="11009" />
                    <RANKING order="4" place="4" resultid="11524" />
                    <RANKING order="5" place="5" resultid="11568" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1307" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11032" />
                    <RANKING order="2" place="2" resultid="11027" />
                    <RANKING order="3" place="3" resultid="11665" />
                    <RANKING order="4" place="-1" resultid="11669" />
                    <RANKING order="5" place="-1" resultid="10979" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11823" daytime="18:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11824" daytime="18:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11825" daytime="18:24" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11826" daytime="18:26" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1308" daytime="18:28" gender="F" number="39" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1309" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11396" />
                    <RANKING order="2" place="2" resultid="11450" />
                    <RANKING order="3" place="3" resultid="10966" />
                    <RANKING order="4" place="4" resultid="11508" />
                    <RANKING order="5" place="-1" resultid="11621" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1310" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11707" />
                    <RANKING order="2" place="2" resultid="10947" />
                    <RANKING order="3" place="3" resultid="10951" />
                    <RANKING order="4" place="4" resultid="11495" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1311" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10853" />
                    <RANKING order="2" place="2" resultid="11702" />
                    <RANKING order="3" place="3" resultid="11419" />
                    <RANKING order="4" place="4" resultid="11633" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1312" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10909" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1313" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10913" />
                    <RANKING order="2" place="2" resultid="10924" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1314" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="11112" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1315" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11101" />
                    <RANKING order="2" place="-1" resultid="11684" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11827" daytime="18:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11828" daytime="18:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11829" daytime="18:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11830" daytime="18:36" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1316" daytime="18:40" gender="M" number="40" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1317" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10975" />
                    <RANKING order="2" place="2" resultid="11455" />
                    <RANKING order="3" place="3" resultid="10987" />
                    <RANKING order="4" place="4" resultid="11629" />
                    <RANKING order="5" place="5" resultid="11018" />
                    <RANKING order="6" place="6" resultid="10893" />
                    <RANKING order="7" place="7" resultid="11650" />
                    <RANKING order="8" place="8" resultid="11578" />
                    <RANKING order="9" place="9" resultid="11654" />
                    <RANKING order="10" place="10" resultid="11573" />
                    <RANKING order="11" place="11" resultid="11645" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1318" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11248" />
                    <RANKING order="2" place="2" resultid="11438" />
                    <RANKING order="3" place="3" resultid="11131" />
                    <RANKING order="4" place="4" resultid="10858" />
                    <RANKING order="5" place="5" resultid="11400" />
                    <RANKING order="6" place="6" resultid="11692" />
                    <RANKING order="7" place="7" resultid="11642" />
                    <RANKING order="8" place="8" resultid="11593" />
                    <RANKING order="9" place="9" resultid="11516" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1319" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10874" />
                    <RANKING order="2" place="2" resultid="11245" />
                    <RANKING order="3" place="3" resultid="10931" />
                    <RANKING order="4" place="4" resultid="11637" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1320" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10869" />
                    <RANKING order="2" place="2" resultid="11610" />
                    <RANKING order="3" place="3" resultid="11598" />
                    <RANKING order="4" place="4" resultid="11662" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1321" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10878" />
                    <RANKING order="2" place="2" resultid="11108" />
                    <RANKING order="3" place="-1" resultid="11443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1322" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11105" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1323" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11233" />
                    <RANKING order="2" place="2" resultid="11602" />
                    <RANKING order="3" place="3" resultid="10954" />
                    <RANKING order="4" place="4" resultid="11615" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11831" daytime="18:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11832" daytime="18:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11833" daytime="18:44" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11834" daytime="18:46" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11835" daytime="18:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="11836" daytime="18:52" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1324" daytime="18:54" gender="F" number="41" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11718" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11157" />
                    <RANKING order="2" place="2" resultid="11162" />
                    <RANKING order="3" place="3" resultid="11172" />
                    <RANKING order="4" place="4" resultid="11182" />
                    <RANKING order="5" place="5" resultid="11152" />
                    <RANKING order="6" place="6" resultid="11147" />
                    <RANKING order="7" place="7" resultid="11545" />
                    <RANKING order="8" place="8" resultid="11207" />
                    <RANKING order="9" place="9" resultid="11202" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11837" daytime="18:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11838" daytime="18:56" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1326" daytime="18:58" gender="M" number="42" order="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11719" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11563" />
                    <RANKING order="2" place="2" resultid="11177" />
                    <RANKING order="3" place="3" resultid="11686" />
                    <RANKING order="4" place="4" resultid="11137" />
                    <RANKING order="5" place="5" resultid="11217" />
                    <RANKING order="6" place="6" resultid="11142" />
                    <RANKING order="7" place="7" resultid="11222" />
                    <RANKING order="8" place="8" resultid="11167" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11839" daytime="18:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11840" daytime="19:02" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1328" daytime="19:04" gender="F" number="43" order="23" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1329" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="1330" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11037" />
                    <RANKING order="2" place="2" resultid="11503" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11841" daytime="19:04" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1331" daytime="19:08" gender="M" number="44" order="24" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1332" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11126" />
                    <RANKING order="2" place="2" resultid="11087" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1333" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11356" />
                    <RANKING order="2" place="2" resultid="11485" />
                    <RANKING order="3" place="3" resultid="11062" />
                    <RANKING order="4" place="4" resultid="11364" />
                    <RANKING order="5" place="5" resultid="11014" />
                    <RANKING order="6" place="6" resultid="11121" />
                    <RANKING order="7" place="7" resultid="11557" />
                    <RANKING order="8" place="8" resultid="11092" />
                    <RANKING order="9" place="-1" resultid="11499" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11842" daytime="19:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11843" daytime="19:10" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1334" daytime="19:14" gender="F" number="45" order="25" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1335" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11328" />
                    <RANKING order="2" place="2" resultid="11082" />
                    <RANKING order="3" place="3" resultid="11000" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1336" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11379" />
                    <RANKING order="2" place="2" resultid="10960" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1337" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11333" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1338" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11337" />
                    <RANKING order="2" place="2" resultid="11496" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1339" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="10848" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1340" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1341" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11230" />
                    <RANKING order="2" place="-1" resultid="11135" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1342" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1343" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11844" daytime="19:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11845" daytime="19:20" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1344" daytime="19:24" gender="M" number="46" order="26" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1345" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11005" />
                    <RANKING order="2" place="2" resultid="11292" />
                    <RANKING order="3" place="3" resultid="11053" />
                    <RANKING order="4" place="4" resultid="11073" />
                    <RANKING order="5" place="5" resultid="11351" />
                    <RANKING order="6" place="6" resultid="11117" />
                    <RANKING order="7" place="7" resultid="11370" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1346" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11323" />
                    <RANKING order="2" place="2" resultid="11282" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1347" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10983" />
                    <RANKING order="2" place="2" resultid="11317" />
                    <RANKING order="3" place="3" resultid="11630" />
                    <RANKING order="4" place="4" resultid="11269" />
                    <RANKING order="5" place="5" resultid="11347" />
                    <RANKING order="6" place="6" resultid="11456" />
                    <RANKING order="7" place="7" resultid="11651" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1348" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11429" />
                    <RANKING order="2" place="2" resultid="11434" />
                    <RANKING order="3" place="3" resultid="11288" />
                    <RANKING order="4" place="-1" resultid="11341" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1349" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11307" />
                    <RANKING order="2" place="2" resultid="11264" />
                    <RANKING order="3" place="3" resultid="11362" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1350" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11612" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1351" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11242" />
                    <RANKING order="2" place="2" resultid="10917" />
                    <RANKING order="3" place="3" resultid="10937" />
                    <RANKING order="4" place="4" resultid="10886" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1352" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="11237" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1353" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="11603" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="11846" daytime="19:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="11847" daytime="19:28" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="11848" daytime="19:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="11849" daytime="19:38" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="11850" daytime="19:40" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="13025" nation="BRA" region="PR" clubid="11226" name="Instituto Desportos Aquáticos De Foz Do Iguaçu" shortname="Cataratas Natação">
          <ATHLETES>
            <ATHLETE firstname="Christopher" lastname="De Araujo" birthdate="2008-08-09" gender="M" nation="BRA" license="366376" athleteid="11238" externalid="366376" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1068" status="DNS" swimtime="00:00:00.00" resultid="11239" heatid="11726" lane="2" entrytime="00:02:00.30" entrycourse="SCM" />
                <RESULT eventid="1094" points="461" swimtime="00:02:35.53" resultid="11240" heatid="11733" lane="2" entrytime="00:02:40.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                    <SPLIT distance="100" swimtime="00:01:13.91" />
                    <SPLIT distance="150" swimtime="00:01:55.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="475" swimtime="00:01:10.80" resultid="11241" heatid="11797" lane="5" entrytime="00:01:12.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="504" swimtime="00:02:17.71" resultid="11242" heatid="11850" lane="4" entrytime="00:02:19.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.28" />
                    <SPLIT distance="100" swimtime="00:01:04.96" />
                    <SPLIT distance="150" swimtime="00:01:45.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Resende Ames" birthdate="2010-02-02" gender="M" nation="BRA" license="365505" athleteid="11250" externalid="365505" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1152" points="352" swimtime="00:01:07.66" resultid="11251" heatid="11757" lane="3" entrytime="00:01:06.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="373" swimtime="00:02:28.40" resultid="11252" heatid="11814" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                    <SPLIT distance="100" swimtime="00:01:07.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Resende Ames" birthdate="2006-02-10" gender="M" nation="BRA" license="365657" athleteid="11234" externalid="365657" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1068" status="DNS" swimtime="00:00:00.00" resultid="11235" heatid="11726" lane="4" entrytime="00:01:58.04" entrycourse="SCM" />
                <RESULT eventid="1270" status="DNS" swimtime="00:00:00.00" resultid="11236" heatid="11810" lane="3" entrytime="00:02:14.84" entrycourse="SCM" />
                <RESULT eventid="1344" status="DNS" swimtime="00:00:00.00" resultid="11237" heatid="11850" lane="3" entrytime="00:02:16.92" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Faisal" lastname="Basem Ghotme" birthdate="2010-12-18" gender="M" nation="BRA" license="390809" athleteid="11243" externalid="390809" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1170" points="502" swimtime="00:00:25.35" resultid="11244" heatid="11767" lane="5" entrytime="00:00:25.98" entrycourse="SCM" />
                <RESULT eventid="1316" points="468" swimtime="00:00:57.73" resultid="11245" heatid="11835" lane="3" entrytime="00:00:58.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Carvalho Carelli" birthdate="2011-10-15" gender="M" nation="BRA" license="403146" athleteid="11246" externalid="403146" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1068" points="457" swimtime="00:02:08.94" resultid="11247" heatid="11726" lane="1" entrytime="00:02:08.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                    <SPLIT distance="100" swimtime="00:01:02.72" />
                    <SPLIT distance="150" swimtime="00:01:35.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="403" swimtime="00:01:00.70" resultid="11248" heatid="11835" lane="4" entrytime="00:01:00.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="384" swimtime="00:02:26.96" resultid="11249" heatid="11814" lane="4" entrytime="00:02:44.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="100" swimtime="00:01:10.97" />
                    <SPLIT distance="150" swimtime="00:01:50.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Victor Oliveira" birthdate="2003-07-16" gender="M" nation="BRA" license="295723" athleteid="11231" externalid="295723" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1152" points="500" swimtime="00:01:00.18" resultid="11232" heatid="11758" lane="3" entrytime="00:00:59.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="508" swimtime="00:00:56.16" resultid="11233" heatid="11836" lane="5" entrytime="00:00:56.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Pinheiro" birthdate="2008-09-04" gender="F" nation="BRA" license="331610" athleteid="11227" externalid="331610">
              <RESULTS>
                <RESULT eventid="1112" points="416" reactiontime="+62" swimtime="00:01:13.49" resultid="11228" heatid="11742" lane="2" entrytime="00:01:14.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1262" points="417" reactiontime="+61" swimtime="00:02:39.14" resultid="11229" heatid="11807" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                    <SPLIT distance="100" swimtime="00:01:17.88" />
                    <SPLIT distance="150" swimtime="00:01:59.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="442" swimtime="00:02:39.96" resultid="11230" heatid="11845" lane="3" entrytime="00:02:38.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                    <SPLIT distance="100" swimtime="00:01:14.56" />
                    <SPLIT distance="150" swimtime="00:02:04.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="11880" points="450" swimtime="00:05:37.88" resultid="11897" heatid="11896" lane="6" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                    <SPLIT distance="100" swimtime="00:01:14.60" />
                    <SPLIT distance="150" swimtime="00:01:59.19" />
                    <SPLIT distance="200" swimtime="00:02:42.12" />
                    <SPLIT distance="250" swimtime="00:03:31.95" />
                    <SPLIT distance="300" swimtime="00:04:22.35" />
                    <SPLIT distance="350" swimtime="00:05:01.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2416" nation="BRA" region="PR" clubid="10865" name="Apan/Maringá">
          <ATHLETES>
            <ATHLETE firstname="Daniel" lastname="Vaneti Mazuti" birthdate="2014-11-29" gender="M" nation="BRA" license="414850" athleteid="11113" externalid="414850">
              <RESULTS>
                <RESULT eventid="1183" status="DNS" swimtime="00:00:00.00" resultid="11114" heatid="11774" lane="5" entrytime="00:00:46.13" entrycourse="SCM" />
                <RESULT eventid="1107" points="115" swimtime="00:00:51.26" resultid="11115" heatid="11738" lane="2" entrytime="00:00:51.55" entrycourse="SCM" />
                <RESULT eventid="1238" points="133" swimtime="00:01:48.18" resultid="11116" heatid="11792" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="137" swimtime="00:03:32.41" resultid="11117" heatid="11846" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.87" />
                    <SPLIT distance="100" swimtime="00:01:43.75" />
                    <SPLIT distance="150" swimtime="00:02:43.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Garcia Cavalcante" birthdate="2008-08-11" gender="M" nation="BRA" license="369676" athleteid="10883" externalid="369676">
              <RESULTS>
                <RESULT eventid="1094" status="DNS" swimtime="00:00:00.00" resultid="10884" heatid="11733" lane="5" entrytime="00:02:40.78" entrycourse="SCM" />
                <RESULT eventid="1270" points="319" reactiontime="+83" swimtime="00:02:34.57" resultid="10885" heatid="11809" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="100" swimtime="00:01:15.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="377" reactiontime="+578" swimtime="00:02:31.74" resultid="10886" heatid="11847" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                    <SPLIT distance="100" swimtime="00:01:16.03" />
                    <SPLIT distance="150" swimtime="00:01:57.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Catarina" lastname="Wendt Jesus" birthdate="2013-07-09" gender="F" nation="BRA" license="393778" athleteid="11044" externalid="393778">
              <RESULTS>
                <RESULT eventid="1142" points="320" swimtime="00:01:18.99" resultid="11045" heatid="11751" lane="3" entrytime="00:01:23.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="413" swimtime="00:00:30.79" resultid="11046" heatid="11772" lane="3" entrytime="00:00:30.48" entrycourse="SCM" />
                <RESULT eventid="1298" points="418" swimtime="00:01:07.18" resultid="11047" heatid="11822" lane="4" entrytime="00:01:09.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="386" swimtime="00:01:25.61" resultid="11048" heatid="11790" lane="1" entrytime="00:01:29.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduarda" lastname="Pastre" birthdate="2017-09-26" gender="F" nation="BRA" license="421910" athleteid="11181" externalid="421910">
              <RESULTS>
                <RESULT eventid="1324" points="44" swimtime="00:01:04.67" resultid="11182" heatid="11838" lane="4" entrytime="00:00:56.97" entrycourse="SCM" />
                <RESULT eventid="1258" points="87" swimtime="00:00:26.77" resultid="11183" heatid="11804" lane="2" entrytime="00:00:27.89" entrycourse="SCM" />
                <RESULT eventid="1224" points="57" swimtime="00:00:34.12" resultid="11184" heatid="11785" lane="1" />
                <RESULT eventid="1294" points="60" swimtime="00:00:28.50" resultid="11185" heatid="11817" lane="4" entrytime="00:00:31.03" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Campos" birthdate="2013-02-17" gender="M" nation="BRA" license="377262" athleteid="10976" externalid="377262">
              <RESULTS>
                <RESULT eventid="1152" status="SICK" swimtime="00:00:00.00" resultid="10977" heatid="11755" lane="6" entrytime="00:01:45.16" entrycourse="SCM" />
                <RESULT eventid="1122" status="SICK" swimtime="00:00:00.00" resultid="10978" heatid="11744" lane="4" entrytime="00:01:27.26" entrycourse="SCM" />
                <RESULT eventid="1303" status="SICK" swimtime="00:00:00.00" resultid="10979" heatid="11826" lane="2" entrytime="00:01:20.16" entrycourse="SCM" />
                <RESULT eventid="1253" status="SICK" swimtime="00:00:00.00" resultid="10980" heatid="11802" lane="4" entrytime="00:00:39.04" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Pedroso Chaim" birthdate="2017-06-14" gender="F" nation="BRA" license="421914" athleteid="11201" externalid="421914">
              <RESULTS>
                <RESULT eventid="1324" points="16" swimtime="00:01:30.18" resultid="11202" heatid="11837" lane="3" />
                <RESULT eventid="1258" points="27" swimtime="00:00:39.20" resultid="11203" heatid="11803" lane="2" />
                <RESULT eventid="1224" points="17" swimtime="00:00:50.78" resultid="11204" heatid="11785" lane="5" entrytime="00:00:52.28" entrycourse="SCM" />
                <RESULT eventid="1294" points="13" swimtime="00:00:46.83" resultid="11205" heatid="11816" lane="2" entrytime="00:00:38.11" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Biason Santana" birthdate="2009-01-21" gender="M" nation="BRA" license="366969" athleteid="10918" externalid="366969">
              <RESULTS>
                <RESULT eventid="1152" points="442" swimtime="00:01:02.69" resultid="10919" heatid="11758" lane="6" entrytime="00:01:02.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="388" swimtime="00:02:26.49" resultid="10920" heatid="11815" lane="5" entrytime="00:02:28.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="100" swimtime="00:01:08.18" />
                    <SPLIT distance="150" swimtime="00:01:46.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Yumi Boso" birthdate="2017-11-26" gender="F" nation="BRA" license="421908" athleteid="11171" externalid="421908">
              <RESULTS>
                <RESULT eventid="1324" points="58" swimtime="00:00:59.15" resultid="11172" heatid="11838" lane="1" />
                <RESULT eventid="1258" points="65" swimtime="00:00:29.50" resultid="11173" heatid="11804" lane="1" entrytime="00:00:30.60" entrycourse="SCM" />
                <RESULT eventid="1224" points="66" swimtime="00:00:32.53" resultid="11174" heatid="11785" lane="3" entrytime="00:00:32.50" entrycourse="SCM" />
                <RESULT eventid="1294" points="39" swimtime="00:00:32.88" resultid="11175" heatid="11817" lane="5" entrytime="00:00:34.03" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raphael" lastname="Piai Pellegrini" birthdate="2012-03-24" gender="M" nation="BRA" license="377261" athleteid="10973" externalid="377261">
              <RESULTS>
                <RESULT eventid="1170" points="415" swimtime="00:00:27.02" resultid="10974" heatid="11766" lane="4" entrytime="00:00:28.37" entrycourse="SCM" />
                <RESULT eventid="1316" points="420" swimtime="00:00:59.83" resultid="10975" heatid="11835" lane="6" entrytime="00:01:03.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathan" lastname="Novak Pinho" birthdate="2012-11-14" gender="M" nation="BRA" license="378199" athleteid="10985" externalid="378199">
              <RESULTS>
                <RESULT eventid="1122" points="219" swimtime="00:01:20.06" resultid="10986" heatid="11744" lane="3" entrytime="00:01:24.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="278" swimtime="00:01:08.63" resultid="10987" heatid="11833" lane="1" entrytime="00:01:17.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Rampasi" birthdate="2013-10-16" gender="F" nation="BRA" license="382209" athleteid="10991" externalid="382209">
              <RESULTS>
                <RESULT eventid="1112" points="133" reactiontime="+79" swimtime="00:01:47.41" resultid="10992" heatid="11739" lane="3" />
                <RESULT eventid="1102" points="154" swimtime="00:00:52.91" resultid="10993" heatid="11736" lane="2" entrytime="00:00:55.26" entrycourse="SCM" />
                <RESULT eventid="1298" points="167" swimtime="00:01:31.14" resultid="10994" heatid="11821" lane="2" entrytime="00:01:26.72" entrycourse="SCM" />
                <RESULT eventid="1204" points="196" swimtime="00:06:37.77" resultid="10995" heatid="11779" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Munhos Donato" birthdate="2016-07-11" gender="F" nation="BRA" license="421912" athleteid="11191" externalid="421912">
              <RESULTS>
                <RESULT eventid="1132" points="36" swimtime="00:01:13.59" resultid="11192" heatid="11747" lane="5" entrytime="00:01:09.94" entrycourse="SCM" />
                <RESULT eventid="1178" points="72" swimtime="00:00:54.88" resultid="11193" heatid="11769" lane="6" entrytime="00:00:54.75" entrycourse="SCM" />
                <RESULT eventid="1298" points="64" swimtime="00:02:05.14" resultid="11194" heatid="11819" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="51" reactiontime="+66" swimtime="00:01:08.01" resultid="11195" heatid="11798" lane="3" entrytime="00:01:04.83" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Pavão" birthdate="2012-04-04" gender="F" nation="BRA" license="377259" athleteid="10964" externalid="377259">
              <RESULTS>
                <RESULT eventid="1112" points="325" reactiontime="+59" swimtime="00:01:19.83" resultid="10965" heatid="11741" lane="2" entrytime="00:01:22.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1308" points="325" swimtime="00:01:13.08" resultid="10966" heatid="11829" lane="1" entrytime="00:01:13.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1262" points="329" reactiontime="+60" swimtime="00:02:52.20" resultid="10967" heatid="11807" lane="3" entrytime="00:02:56.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.83" />
                    <SPLIT distance="100" swimtime="00:01:24.18" />
                    <SPLIT distance="150" swimtime="00:02:08.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio" lastname="Rafael Padial" birthdate="2014-03-07" gender="M" nation="BRA" license="397331" athleteid="11049" externalid="397331">
              <RESULTS>
                <RESULT eventid="1122" points="144" swimtime="00:01:32.12" resultid="11050" heatid="11744" lane="5" entrytime="00:01:35.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="180" swimtime="00:00:35.65" resultid="11051" heatid="11776" lane="1" entrytime="00:00:35.06" entrycourse="SCM" />
                <RESULT eventid="1303" points="182" swimtime="00:01:19.01" resultid="11052" heatid="11826" lane="5" entrytime="00:01:20.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="163" swimtime="00:03:20.60" resultid="11053" heatid="11847" lane="4" entrytime="00:03:26.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Peroni Passafaro" birthdate="2013-09-17" gender="F" nation="BRA" license="370659" athleteid="10956" externalid="370659">
              <RESULTS>
                <RESULT eventid="1112" points="277" reactiontime="+76" swimtime="00:01:24.18" resultid="10957" heatid="11740" lane="4" entrytime="00:01:27.64" entrycourse="SCM" />
                <RESULT eventid="1178" points="318" swimtime="00:00:33.56" resultid="10958" heatid="11772" lane="6" entrytime="00:00:35.21" entrycourse="SCM" />
                <RESULT comment="SW 7.1 - Mais de uma pernada de borboleta antes da primeira pernada de peito após o início ou a virada., Na volta dos 25m." eventid="1228" status="DSQ" swimtime="00:01:48.85" resultid="10959" heatid="11789" lane="5" entrytime="00:01:56.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="253" swimtime="00:03:12.56" resultid="10960" heatid="11845" lane="6" entrytime="00:03:25.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.11" />
                    <SPLIT distance="100" swimtime="00:01:31.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lavinia" lastname="Bossoni" birthdate="2013-11-03" gender="F" nation="BRA" license="377260" athleteid="10968" externalid="377260">
              <RESULTS>
                <RESULT eventid="1112" points="181" reactiontime="+67" swimtime="00:01:37.02" resultid="10969" heatid="11740" lane="1" entrytime="00:01:38.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="263" swimtime="00:00:35.76" resultid="10970" heatid="11771" lane="2" entrytime="00:00:39.07" entrycourse="SCM" />
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Tempo: 16:38), Na volta dos 25m." eventid="1228" status="DSQ" swimtime="00:01:47.01" resultid="10971" heatid="11789" lane="2" entrytime="00:01:46.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="190" swimtime="00:06:42.20" resultid="10972" heatid="11779" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.38" />
                    <SPLIT distance="100" swimtime="00:01:38.62" />
                    <SPLIT distance="150" swimtime="00:02:31.38" />
                    <SPLIT distance="200" swimtime="00:03:23.01" />
                    <SPLIT distance="250" swimtime="00:04:14.82" />
                    <SPLIT distance="300" swimtime="00:05:04.86" />
                    <SPLIT distance="350" swimtime="00:05:55.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Marques Picolo Vinha" birthdate="2010-07-01" gender="M" nation="BRA" license="366990" athleteid="10929" externalid="366990">
              <RESULTS>
                <RESULT eventid="1170" points="370" swimtime="00:00:28.07" resultid="10930" heatid="11766" lane="2" entrytime="00:00:28.48" entrycourse="SCM" />
                <RESULT eventid="1316" points="384" swimtime="00:01:01.69" resultid="10931" heatid="11834" lane="3" entrytime="00:01:03.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Sanches Ghelere" birthdate="2008-08-06" gender="F" nation="BRA" license="372024" athleteid="10910" externalid="372024">
              <RESULTS>
                <RESULT eventid="1142" points="411" swimtime="00:01:12.69" resultid="10911" heatid="11752" lane="2" entrytime="00:01:16.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="506" swimtime="00:02:18.40" resultid="10912" heatid="11723" lane="1" entrytime="00:02:25.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                    <SPLIT distance="100" swimtime="00:01:06.35" />
                    <SPLIT distance="150" swimtime="00:01:42.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1308" points="520" swimtime="00:01:02.45" resultid="10913" heatid="11830" lane="4" entrytime="00:01:02.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edgar" lastname="Romero" birthdate="2011-05-12" gender="M" nation="BRA" license="413920" athleteid="11128" externalid="413920">
              <RESULTS>
                <RESULT eventid="1068" points="275" swimtime="00:02:32.68" resultid="11129" heatid="11724" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.45" />
                    <SPLIT distance="100" swimtime="00:01:11.51" />
                    <SPLIT distance="150" swimtime="00:01:53.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="314" swimtime="00:00:29.63" resultid="11130" heatid="11764" lane="4" entrytime="00:00:32.74" entrycourse="SCM" />
                <RESULT eventid="1316" points="314" swimtime="00:01:05.93" resultid="11131" heatid="11834" lane="6" entrytime="00:01:12.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Antonio Mendes" birthdate="2008-12-04" gender="M" nation="BRA" license="366962" athleteid="10914" externalid="366962">
              <RESULTS>
                <RESULT eventid="1122" points="437" swimtime="00:01:03.68" resultid="10915" heatid="11874" lane="3" entrytime="00:01:04.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="413" reactiontime="+63" swimtime="00:02:21.79" resultid="10916" heatid="11810" lane="4" entrytime="00:02:19.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                    <SPLIT distance="100" swimtime="00:01:07.52" />
                    <SPLIT distance="150" swimtime="00:01:44.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="495" swimtime="00:02:18.53" resultid="10917" heatid="11850" lane="2" entrytime="00:02:23.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juan" lastname="Bernardo Padua" birthdate="2013-07-15" gender="M" nation="BRA" license="392108" athleteid="11019" externalid="392108">
              <RESULTS>
                <RESULT eventid="1183" points="224" swimtime="00:00:33.19" resultid="11020" heatid="11776" lane="5" entrytime="00:00:34.66" entrycourse="SCM" />
                <RESULT eventid="1137" points="206" swimtime="00:00:36.79" resultid="11021" heatid="11749" lane="4" entrytime="00:00:38.33" entrycourse="SCM" />
                <RESULT eventid="1238" points="184" swimtime="00:01:37.14" resultid="11022" heatid="11794" lane="4" entrytime="00:01:37.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1214" points="200" swimtime="00:06:02.79" resultid="11023" heatid="11782" lane="1" entrytime="00:06:11.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                    <SPLIT distance="100" swimtime="00:01:27.30" />
                    <SPLIT distance="150" swimtime="00:02:13.96" />
                    <SPLIT distance="200" swimtime="00:03:00.40" />
                    <SPLIT distance="250" swimtime="00:03:47.40" />
                    <SPLIT distance="300" swimtime="00:04:34.61" />
                    <SPLIT distance="350" swimtime="00:05:21.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Cristina Mussolim" birthdate="2015-05-16" gender="F" nation="BRA" license="421913" athleteid="11196" externalid="421913">
              <RESULTS>
                <RESULT eventid="1178" points="107" swimtime="00:00:48.17" resultid="11197" heatid="11769" lane="4" entrytime="00:00:50.50" entrycourse="SCM" />
                <RESULT eventid="1102" points="64" swimtime="00:01:10.67" resultid="11198" heatid="11735" lane="1" entrytime="00:01:07.23" entrycourse="SCM" />
                <RESULT eventid="1298" points="101" swimtime="00:01:47.69" resultid="11199" heatid="11819" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="81" reactiontime="+95" swimtime="00:00:58.33" resultid="11200" heatid="11799" lane="1" entrytime="00:01:03.44" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Casavechia Carraro" birthdate="2009-07-28" gender="M" nation="BRA" license="368150" athleteid="10866" externalid="368150">
              <RESULTS>
                <RESULT eventid="1068" points="646" swimtime="00:01:54.91" resultid="10867" heatid="11726" lane="3" entrytime="00:01:55.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.98" />
                    <SPLIT distance="100" swimtime="00:00:56.74" />
                    <SPLIT distance="150" swimtime="00:01:25.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="483" swimtime="00:00:25.69" resultid="10868" heatid="11767" lane="3" entrytime="00:00:24.72" entrycourse="SCM" />
                <RESULT eventid="1316" points="653" swimtime="00:00:51.66" resultid="10869" heatid="11836" lane="3" entrytime="00:00:51.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="489" swimtime="00:02:15.60" resultid="10870" heatid="11813" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.31" />
                    <SPLIT distance="100" swimtime="00:01:03.40" />
                    <SPLIT distance="150" swimtime="00:01:38.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heitor" lastname="Bello Paula" birthdate="2015-06-14" gender="M" nation="BRA" license="393776" athleteid="11039" externalid="393776">
              <RESULTS>
                <RESULT eventid="1183" points="125" swimtime="00:00:40.32" resultid="11040" heatid="11775" lane="1" entrytime="00:00:39.35" entrycourse="SCM" />
                <RESULT eventid="1107" points="90" reactiontime="+198" swimtime="00:00:55.64" resultid="11041" heatid="11738" lane="1" entrytime="00:00:55.85" entrycourse="SCM" />
                <RESULT eventid="1303" points="103" swimtime="00:01:35.42" resultid="11042" heatid="11825" lane="6" entrytime="00:01:37.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1253" points="91" reactiontime="+79" swimtime="00:00:49.09" resultid="11043" heatid="11802" lane="6" entrytime="00:00:46.58" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniela" lastname="Inoue" birthdate="2008-10-31" gender="F" nation="BRA" license="378348" athleteid="10921" externalid="378348">
              <RESULTS>
                <RESULT eventid="1112" points="269" reactiontime="+71" swimtime="00:01:24.94" resultid="10922" heatid="11741" lane="1" entrytime="00:01:23.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1162" points="373" swimtime="00:00:31.83" resultid="10923" heatid="11761" lane="5" entrytime="00:00:31.33" entrycourse="SCM" />
                <RESULT eventid="1308" points="350" swimtime="00:01:11.24" resultid="10924" heatid="11829" lane="4" entrytime="00:01:10.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Da Cateburcio" birthdate="2004-01-18" gender="F" nation="BRA" license="407186" athleteid="11099" externalid="407186">
              <RESULTS>
                <RESULT eventid="1162" points="96" swimtime="00:00:50.03" resultid="11100" heatid="11759" lane="5" entrytime="00:00:52.12" entrycourse="SCM" />
                <RESULT eventid="1308" points="92" swimtime="00:01:50.95" resultid="11101" heatid="11827" lane="4" entrytime="00:01:58.78" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Dos Reis Monteiro" birthdate="2014-08-05" gender="M" nation="BRA" license="392095" athleteid="11001" externalid="392095">
              <RESULTS>
                <RESULT eventid="1152" points="179" swimtime="00:01:24.70" resultid="11002" heatid="11753" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="231" swimtime="00:00:32.83" resultid="11003" heatid="11776" lane="3" entrytime="00:00:32.22" entrycourse="SCM" />
                <RESULT eventid="1238" points="227" swimtime="00:01:30.59" resultid="11004" heatid="11795" lane="6" entrytime="00:01:35.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="224" swimtime="00:03:00.37" resultid="11005" heatid="11848" lane="6" entrytime="00:03:06.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                    <SPLIT distance="100" swimtime="00:01:30.06" />
                    <SPLIT distance="150" swimtime="00:02:19.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Izzo Campos" birthdate="2017-05-29" gender="M" nation="BRA" license="421960" athleteid="11216" externalid="421960">
              <RESULTS>
                <RESULT eventid="1326" points="42" swimtime="00:00:57.56" resultid="11217" heatid="11840" lane="3" entrytime="00:00:54.74" entrycourse="SCM" />
                <RESULT eventid="1226" points="41" swimtime="00:00:33.17" resultid="11218" heatid="11786" lane="3" />
                <RESULT eventid="1260" points="35" swimtime="00:00:31.38" resultid="11219" heatid="11806" lane="4" entrytime="00:00:29.99" entrycourse="SCM" />
                <RESULT eventid="1296" points="25" swimtime="00:00:33.56" resultid="11220" heatid="11818" lane="5" entrytime="00:00:33.33" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carina" lastname="Costa Profeta" birthdate="2008-03-20" gender="F" nation="BRA" license="366964" athleteid="10904" externalid="366964">
              <RESULTS>
                <RESULT eventid="1162" points="435" swimtime="00:00:30.26" resultid="10905" heatid="11761" lane="4" entrytime="00:00:30.78" entrycourse="SCM" />
                <RESULT eventid="1228" points="447" swimtime="00:01:21.55" resultid="10906" heatid="11791" lane="5" entrytime="00:01:19.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Marques" birthdate="2015-10-15" gender="F" nation="BRA" license="399738" athleteid="11064" externalid="399738">
              <RESULTS>
                <RESULT eventid="1132" points="47" swimtime="00:01:07.35" resultid="11065" heatid="11747" lane="1" entrytime="00:01:29.26" entrycourse="SCM" />
                <RESULT eventid="1178" points="89" swimtime="00:00:51.34" resultid="11066" heatid="11768" lane="3" entrytime="00:00:55.51" entrycourse="SCM" />
                <RESULT eventid="1298" points="68" swimtime="00:02:02.53" resultid="11067" heatid="11820" lane="4" entrytime="00:02:00.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="67" reactiontime="+69" swimtime="00:01:02.11" resultid="11068" heatid="11799" lane="5" entrytime="00:01:01.40" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Ayres" birthdate="2012-05-05" gender="M" nation="BRA" license="378035" athleteid="10981" externalid="378035">
              <RESULTS>
                <RESULT eventid="1122" points="300" swimtime="00:01:12.14" resultid="10982" heatid="11746" lane="1" entrytime="00:01:12.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="324" swimtime="00:02:39.54" resultid="10983" heatid="11849" lane="5" entrytime="00:02:43.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.71" />
                    <SPLIT distance="100" swimtime="00:01:15.70" />
                    <SPLIT distance="150" swimtime="00:02:04.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1214" points="362" swimtime="00:04:57.63" resultid="10984" heatid="11783" lane="1" entrytime="00:05:00.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.80" />
                    <SPLIT distance="100" swimtime="00:01:10.57" />
                    <SPLIT distance="150" swimtime="00:01:49.45" />
                    <SPLIT distance="200" swimtime="00:02:27.80" />
                    <SPLIT distance="250" swimtime="00:03:05.64" />
                    <SPLIT distance="300" swimtime="00:03:44.60" />
                    <SPLIT distance="350" swimtime="00:04:23.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Lopes Ferreira" birthdate="2008-12-03" gender="F" nation="ESP" license="383455" athleteid="11132" externalid="383455">
              <RESULTS>
                <RESULT eventid="1112" points="286" reactiontime="+68" swimtime="00:01:23.30" resultid="11133" heatid="11741" lane="6" entrytime="00:01:26.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1162" points="275" swimtime="00:00:35.25" resultid="11134" heatid="11759" lane="3" entrytime="00:00:37.82" entrycourse="SCM" />
                <RESULT comment="SW 6.2 - Deixou a posição de costas, exceto ao executar uma virada.  (Tempo: 19:31), Costas, Medley Individual." eventid="1334" status="DSQ" swimtime="00:03:18.18" resultid="11135" heatid="11844" lane="1">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:02:36.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Muniz" birthdate="2012-09-03" gender="M" nation="BRA" license="392106" athleteid="11016" externalid="392106">
              <RESULTS>
                <RESULT eventid="1170" points="265" swimtime="00:00:31.35" resultid="11017" heatid="11764" lane="5" entrytime="00:00:33.14" entrycourse="SCM" />
                <RESULT eventid="1316" points="263" swimtime="00:01:09.93" resultid="11018" heatid="11833" lane="3" entrytime="00:01:13.68" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Amelia Sales" birthdate="2017-07-05" gender="F" nation="BRA" license="421906" athleteid="11161" externalid="421906">
              <RESULTS>
                <RESULT eventid="1324" points="61" swimtime="00:00:58.09" resultid="11162" heatid="11838" lane="2" entrytime="00:00:58.01" entrycourse="SCM" />
                <RESULT eventid="1258" points="101" swimtime="00:00:25.42" resultid="11163" heatid="11804" lane="4" entrytime="00:00:26.77" entrycourse="SCM" />
                <RESULT eventid="1224" points="47" swimtime="00:00:36.52" resultid="11164" heatid="11784" lane="4" />
                <RESULT eventid="1294" points="59" swimtime="00:00:28.72" resultid="11165" heatid="11817" lane="2" entrytime="00:00:32.28" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Henrique Goes" birthdate="2008-10-26" gender="M" nation="BRA" license="392105" athleteid="10925" externalid="392105">
              <RESULTS>
                <RESULT eventid="1068" points="304" swimtime="00:02:27.65" resultid="10926" heatid="11725" lane="6" entrytime="00:02:24.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                    <SPLIT distance="100" swimtime="00:01:09.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="248" swimtime="00:01:27.98" resultid="10927" heatid="11795" lane="3" entrytime="00:01:28.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1214" points="266" swimtime="00:05:29.89" resultid="10928" heatid="11782" lane="2" entrytime="00:05:22.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                    <SPLIT distance="100" swimtime="00:01:16.84" />
                    <SPLIT distance="150" swimtime="00:01:58.59" />
                    <SPLIT distance="200" swimtime="00:02:40.75" />
                    <SPLIT distance="250" swimtime="00:03:22.98" />
                    <SPLIT distance="300" swimtime="00:04:05.02" />
                    <SPLIT distance="350" swimtime="00:04:47.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Beffa Silva" birthdate="2017-02-19" gender="M" nation="BRA" license="421902" athleteid="11141" externalid="421902">
              <RESULTS>
                <RESULT eventid="1326" points="34" swimtime="00:01:01.89" resultid="11142" heatid="11840" lane="5" entrytime="00:01:02.85" entrycourse="SCM" />
                <RESULT eventid="1226" points="60" swimtime="00:00:29.24" resultid="11143" heatid="11787" lane="4" entrytime="00:00:37.53" entrycourse="SCM" />
                <RESULT eventid="1260" points="32" swimtime="00:00:32.14" resultid="11144" heatid="11805" lane="3" />
                <RESULT eventid="1296" points="27" swimtime="00:00:32.62" resultid="11145" heatid="11818" lane="4" entrytime="00:00:32.85" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Diogo" lastname="Sanchez" birthdate="2012-11-29" gender="M" nation="BRA" license="370658" athleteid="10890" externalid="370658">
              <RESULTS>
                <RESULT eventid="1094" points="203" swimtime="00:03:24.36" resultid="10891" heatid="11732" lane="5" entrytime="00:03:40.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="211" swimtime="00:00:33.83" resultid="10892" heatid="11763" lane="3" entrytime="00:00:36.70" entrycourse="SCM" />
                <RESULT eventid="1316" points="187" swimtime="00:01:18.36" resultid="10893" heatid="11833" lane="6" entrytime="00:01:19.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="206" swimtime="00:01:33.60" resultid="10894" heatid="11795" lane="2" entrytime="00:01:32.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Chaim" birthdate="2011-05-29" gender="F" nation="BRA" license="370662" athleteid="10945" externalid="370662">
              <RESULTS>
                <RESULT eventid="1162" points="346" swimtime="00:00:32.64" resultid="10946" heatid="11760" lane="4" entrytime="00:00:32.45" entrycourse="SCM" />
                <RESULT eventid="1308" points="345" swimtime="00:01:11.60" resultid="10947" heatid="11829" lane="5" entrytime="00:01:11.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Fernanda Silva Simoes" birthdate="2017-09-05" gender="F" nation="BRA" license="421904" athleteid="11151" externalid="421904">
              <RESULTS>
                <RESULT eventid="1324" points="40" swimtime="00:01:06.50" resultid="11152" heatid="11838" lane="5" entrytime="00:01:09.33" entrycourse="SCM" />
                <RESULT eventid="1258" points="54" swimtime="00:00:31.33" resultid="11153" heatid="11804" lane="5" entrytime="00:00:30.56" entrycourse="SCM" />
                <RESULT eventid="1224" points="46" swimtime="00:00:36.56" resultid="11154" heatid="11785" lane="6" />
                <RESULT eventid="1294" points="29" swimtime="00:00:36.05" resultid="11155" heatid="11817" lane="1" entrytime="00:00:35.15" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio" lastname="Bertalia Souza" birthdate="2017-02-13" gender="M" nation="BRA" license="424506" athleteid="11221" externalid="424506">
              <RESULTS>
                <RESULT eventid="1326" points="34" swimtime="00:01:02.18" resultid="11222" heatid="11839" lane="3" />
                <RESULT eventid="1226" points="59" swimtime="00:00:29.31" resultid="11223" heatid="11786" lane="5" />
                <RESULT eventid="1260" points="28" swimtime="00:00:33.73" resultid="11224" heatid="11806" lane="5" />
                <RESULT eventid="1296" points="27" swimtime="00:00:32.89" resultid="11225" heatid="11818" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Sunahara Machado" birthdate="2015-03-23" gender="M" nation="BRA" license="421911" athleteid="11186" externalid="421911">
              <RESULTS>
                <RESULT eventid="1183" points="52" swimtime="00:00:53.76" resultid="11187" heatid="11773" lane="3" entrytime="00:01:03.67" entrycourse="SCM" />
                <RESULT eventid="1107" points="71" swimtime="00:01:00.09" resultid="11188" heatid="11737" lane="2" entrytime="00:01:05.99" entrycourse="SCM" />
                <RESULT eventid="1303" points="61" swimtime="00:01:53.84" resultid="11189" heatid="11824" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1253" points="30" reactiontime="+80" swimtime="00:01:10.71" resultid="11190" heatid="11801" lane="1" entrytime="00:01:09.37" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Passafaro" birthdate="2009-02-01" gender="F" nation="BRA" license="370673" athleteid="10907" externalid="370673">
              <RESULTS>
                <RESULT eventid="1142" points="317" swimtime="00:01:19.25" resultid="10908" heatid="11752" lane="1" entrytime="00:01:22.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1308" points="343" swimtime="00:01:11.75" resultid="10909" heatid="11830" lane="6" entrytime="00:01:09.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Quental De Meireles" birthdate="2008-11-20" gender="M" nation="BRA" license="392103" athleteid="10935" externalid="392103">
              <RESULTS>
                <RESULT eventid="1152" points="381" swimtime="00:01:05.88" resultid="10936" heatid="11757" lane="2" entrytime="00:01:07.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="378" swimtime="00:02:31.52" resultid="10937" heatid="11846" lane="4">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:01:13.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1214" points="410" swimtime="00:04:45.61" resultid="10938" heatid="11781" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                    <SPLIT distance="100" swimtime="00:01:06.63" />
                    <SPLIT distance="150" swimtime="00:01:42.55" />
                    <SPLIT distance="200" swimtime="00:02:19.78" />
                    <SPLIT distance="250" swimtime="00:02:57.67" />
                    <SPLIT distance="300" swimtime="00:03:35.12" />
                    <SPLIT distance="350" swimtime="00:04:11.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Izzo Breschiliare" birthdate="2015-09-23" gender="M" nation="BRA" license="407182" athleteid="11089" externalid="407182">
              <RESULTS>
                <RESULT eventid="1183" points="109" swimtime="00:00:42.14" resultid="11090" heatid="11774" lane="6" entrytime="00:00:49.73" entrycourse="SCM" />
                <RESULT eventid="1137" points="58" swimtime="00:00:55.92" resultid="11091" heatid="11748" lane="3" entrytime="00:00:58.79" entrycourse="SCM" />
                <RESULT eventid="1331" points="67" swimtime="00:02:00.94" resultid="11092" heatid="11842" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1253" points="72" reactiontime="+65" swimtime="00:00:53.11" resultid="11093" heatid="11801" lane="5" entrytime="00:00:56.67" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Batista Sanchez" birthdate="2009-05-22" gender="M" nation="BRA" license="370668" athleteid="10880" externalid="370668">
              <RESULTS>
                <RESULT eventid="1094" points="383" swimtime="00:02:45.35" resultid="10881" heatid="11733" lane="1" entrytime="00:02:41.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                    <SPLIT distance="100" swimtime="00:01:19.59" />
                    <SPLIT distance="150" swimtime="00:02:02.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="397" swimtime="00:01:15.19" resultid="10882" heatid="11797" lane="2" entrytime="00:01:11.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Bissoli Lucas" birthdate="2017-06-06" gender="M" nation="BRA" license="421907" athleteid="11166" externalid="421907">
              <RESULTS>
                <RESULT eventid="1326" points="30" swimtime="00:01:04.74" resultid="11167" heatid="11840" lane="1" entrytime="00:01:15.61" entrycourse="SCM" />
                <RESULT eventid="1226" points="37" swimtime="00:00:34.23" resultid="11168" heatid="11787" lane="3" entrytime="00:00:36.24" entrycourse="SCM" />
                <RESULT eventid="1260" points="43" swimtime="00:00:29.20" resultid="11169" heatid="11805" lane="2" />
                <RESULT eventid="1296" points="18" swimtime="00:00:37.16" resultid="11170" heatid="11818" lane="1" entrytime="00:00:37.94" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aaron" lastname="Michels Dias" birthdate="2017-07-04" gender="M" nation="BRA" license="421909" athleteid="11176" externalid="421909">
              <RESULTS>
                <RESULT eventid="1326" points="77" swimtime="00:00:47.36" resultid="11177" heatid="11840" lane="4" entrytime="00:00:55.36" entrycourse="SCM" />
                <RESULT eventid="1226" points="59" swimtime="00:00:29.40" resultid="11178" heatid="11786" lane="4" />
                <RESULT eventid="1260" points="86" swimtime="00:00:23.32" resultid="11179" heatid="11806" lane="3" entrytime="00:00:26.10" entrycourse="SCM" />
                <RESULT eventid="1296" points="41" swimtime="00:00:28.41" resultid="11180" heatid="11818" lane="3" entrytime="00:00:27.73" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Fernandes Rivadavia" birthdate="2015-11-15" gender="F" nation="BRA" license="393774" athleteid="11034" externalid="393774">
              <RESULTS>
                <RESULT eventid="1076" points="236" swimtime="00:02:58.40" resultid="11035" heatid="11727" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.62" />
                    <SPLIT distance="100" swimtime="00:01:25.03" />
                    <SPLIT distance="150" swimtime="00:02:13.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="144" swimtime="00:00:46.49" resultid="11036" heatid="11747" lane="2" entrytime="00:00:44.13" entrycourse="SCM" />
                <RESULT eventid="1328" points="215" swimtime="00:01:34.24" resultid="11037" heatid="11841" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="243" swimtime="00:01:20.43" resultid="11038" heatid="11821" lane="4" entrytime="00:01:23.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Isabel Henriques" birthdate="2007-09-05" gender="F" nation="BRA" license="414491" athleteid="11110" externalid="414491">
              <RESULTS>
                <RESULT eventid="1162" status="DNS" swimtime="00:00:00.00" resultid="11111" heatid="11759" lane="4" entrytime="00:00:38.79" entrycourse="SCM" />
                <RESULT eventid="1308" status="DNS" swimtime="00:00:00.00" resultid="11112" heatid="11828" lane="5" entrytime="00:01:29.90" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lara" lastname="Constantino" birthdate="2012-06-02" gender="F" nation="BRA" license="382208" athleteid="10988" externalid="382208">
              <RESULTS>
                <RESULT eventid="1086" points="327" reactiontime="+209" swimtime="00:03:15.20" resultid="10989" heatid="11730" lane="3" entrytime="00:03:25.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.83" />
                    <SPLIT distance="100" swimtime="00:01:35.74" />
                    <SPLIT distance="150" swimtime="00:02:26.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="362" swimtime="00:01:27.47" resultid="10990" heatid="11790" lane="5" entrytime="00:01:29.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Pacheco" birthdate="2012-10-03" gender="M" nation="BRA" license="370663" athleteid="10961" externalid="370663">
              <RESULTS>
                <RESULT eventid="1170" points="287" swimtime="00:00:30.54" resultid="10962" heatid="11765" lane="5" entrytime="00:00:31.27" entrycourse="SCM" />
                <RESULT eventid="1238" points="307" swimtime="00:01:21.88" resultid="10963" heatid="11795" lane="5" entrytime="00:01:33.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Ghelere" birthdate="2011-04-03" gender="F" nation="BRA" license="368146" athleteid="10948" externalid="368146">
              <RESULTS>
                <RESULT eventid="1112" points="344" reactiontime="+76" swimtime="00:01:18.29" resultid="10949" heatid="11741" lane="3" entrytime="00:01:21.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1162" points="330" swimtime="00:00:33.16" resultid="10950" heatid="11760" lane="3" entrytime="00:00:32.30" entrycourse="SCM" />
                <RESULT eventid="1308" points="332" swimtime="00:01:12.53" resultid="10951" heatid="11829" lane="2" entrytime="00:01:10.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tiago" lastname="Ficher Delmont Pais" birthdate="2010-07-15" gender="M" nation="BRA" license="338533" athleteid="10871" externalid="338533">
              <RESULTS>
                <RESULT eventid="1152" points="512" swimtime="00:00:59.71" resultid="10872" heatid="11758" lane="4" entrytime="00:01:00.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="522" swimtime="00:02:03.37" resultid="10873" heatid="11724" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.92" />
                    <SPLIT distance="100" swimtime="00:00:59.06" />
                    <SPLIT distance="150" swimtime="00:01:31.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="521" swimtime="00:00:55.71" resultid="10874" heatid="11836" lane="4" entrytime="00:00:55.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="444" swimtime="00:02:19.96" resultid="10875" heatid="11815" lane="1" entrytime="00:02:33.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.94" />
                    <SPLIT distance="100" swimtime="00:01:04.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Allana" lastname="Araujo Oliveira" birthdate="2017-07-25" gender="F" nation="BRA" license="421905" athleteid="11156" externalid="421905">
              <RESULTS>
                <RESULT eventid="1324" points="97" swimtime="00:00:49.89" resultid="11157" heatid="11838" lane="3" entrytime="00:00:55.40" entrycourse="SCM" />
                <RESULT eventid="1258" points="120" swimtime="00:00:24.05" resultid="11158" heatid="11804" lane="3" entrytime="00:00:23.54" entrycourse="SCM" />
                <RESULT eventid="1224" points="36" swimtime="00:00:39.60" resultid="11159" heatid="11784" lane="3" />
                <RESULT eventid="1294" points="85" swimtime="00:00:25.41" resultid="11160" heatid="11817" lane="3" entrytime="00:00:25.80" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Guilherme Ortega" birthdate="1999-08-05" gender="M" nation="BRA" license="383118" athleteid="10952" externalid="383118">
              <RESULTS>
                <RESULT eventid="1122" points="341" swimtime="00:01:09.17" resultid="10953" heatid="11746" lane="5" entrytime="00:01:09.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="389" swimtime="00:01:01.42" resultid="10954" heatid="11831" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="352" reactiontime="+75" swimtime="00:02:29.54" resultid="10955" heatid="11810" lane="5" entrytime="00:02:35.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                    <SPLIT distance="100" swimtime="00:01:12.90" />
                    <SPLIT distance="150" swimtime="00:01:51.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Tomazeli" birthdate="2013-02-05" gender="M" nation="BRA" license="392109" athleteid="11024" externalid="392109">
              <RESULTS>
                <RESULT comment="SW 8.5 - Totalmente submerso durante o nado.  (Tempo: 11:21)" eventid="1152" status="DSQ" swimtime="00:01:40.37" resultid="11025" heatid="11755" lane="1" entrytime="00:01:42.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="222" swimtime="00:00:33.29" resultid="11026" heatid="11776" lane="4" entrytime="00:00:33.07" entrycourse="SCM" />
                <RESULT eventid="1303" points="191" swimtime="00:01:17.74" resultid="11027" heatid="11823" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="142" swimtime="00:01:45.94" resultid="11028" heatid="11792" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Felipe Sakaguti" birthdate="2007-06-22" gender="M" nation="BRA" license="407187" athleteid="11102" externalid="407187">
              <RESULTS>
                <RESULT eventid="1122" points="96" reactiontime="+112" swimtime="00:01:45.35" resultid="11103" heatid="11743" lane="3" entrytime="00:01:56.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.61" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Tempo: 11:39)" eventid="1170" status="DSQ" swimtime="00:00:40.75" resultid="11104" heatid="11763" lane="1" entrytime="00:00:39.16" entrycourse="SCM" />
                <RESULT eventid="1316" points="113" swimtime="00:01:32.74" resultid="11105" heatid="11832" lane="1" entrytime="00:01:29.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Pastre" birthdate="2014-03-10" gender="F" nation="BRA" license="403760" athleteid="11079" externalid="403760">
              <RESULTS>
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Tempo: 11:06), Na volta dos 25m." eventid="1142" status="DSQ" swimtime="00:01:38.14" resultid="11080" heatid="11750" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="249" reactiontime="+66" swimtime="00:01:27.14" resultid="11081" heatid="11740" lane="5" entrytime="00:01:34.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="220" swimtime="00:03:21.78" resultid="11082" heatid="11844" lane="2" entrytime="00:03:36.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.28" />
                    <SPLIT distance="100" swimtime="00:01:39.02" />
                    <SPLIT distance="150" swimtime="00:02:38.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="279" reactiontime="+68" swimtime="00:00:38.61" resultid="11083" heatid="11800" lane="4" entrytime="00:00:40.03" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Borges Carneiro" birthdate="1998-05-07" gender="F" nation="BRA" license="266382" athleteid="10898" externalid="266382" level="S14 - SM14">
              <RESULTS>
                <RESULT eventid="1086" points="514" status="EXH" swimtime="00:02:47.90" resultid="10899" heatid="11731" lane="4" entrytime="00:02:50.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                    <SPLIT distance="100" swimtime="00:01:18.96" />
                    <SPLIT distance="150" swimtime="00:02:02.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="527" status="EXH" swimtime="00:01:17.16" resultid="10900" heatid="11791" lane="2" entrytime="00:01:18.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="De Araujo" birthdate="2015-08-09" gender="F" nation="BRA" license="407185" athleteid="11094" externalid="407185">
              <RESULTS>
                <RESULT eventid="1178" points="86" swimtime="00:00:51.91" resultid="11095" heatid="11769" lane="1" entrytime="00:00:52.01" entrycourse="SCM" />
                <RESULT eventid="1102" points="98" swimtime="00:01:01.46" resultid="11096" heatid="11736" lane="6" entrytime="00:00:57.79" entrycourse="SCM" />
                <RESULT eventid="1298" points="67" swimtime="00:02:03.70" resultid="11097" heatid="11819" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="63" reactiontime="+113" swimtime="00:01:03.30" resultid="11098" heatid="11799" lane="2" entrytime="00:00:59.09" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hammon" lastname="Henrique Costa" birthdate="2008-09-19" gender="M" nation="BRA" license="408703" athleteid="11106" externalid="408703">
              <RESULTS>
                <RESULT eventid="1170" points="363" swimtime="00:00:28.24" resultid="11107" heatid="11766" lane="3" entrytime="00:00:28.04" entrycourse="SCM" />
                <RESULT eventid="1316" points="318" swimtime="00:01:05.67" resultid="11108" heatid="11834" lane="4" entrytime="00:01:04.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="341" swimtime="00:01:19.07" resultid="11109" heatid="11796" lane="3" entrytime="00:01:18.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Santos Carraro" birthdate="2014-06-04" gender="M" nation="BRA" license="392097" athleteid="11006" externalid="392097">
              <RESULTS>
                <RESULT eventid="1152" points="108" swimtime="00:01:40.08" resultid="11007" heatid="11753" lane="4" />
                <RESULT eventid="1122" points="120" reactiontime="+71" swimtime="00:01:37.94" resultid="11008" heatid="11743" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="164" swimtime="00:01:21.84" resultid="11009" heatid="11826" lane="1" entrytime="00:01:21.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="113" swimtime="00:01:54.26" resultid="11010" heatid="11793" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laion" lastname="Miguel Simoes" birthdate="2016-04-02" gender="M" nation="BRA" license="407179" athleteid="11084" externalid="407179">
              <RESULTS>
                <RESULT eventid="1081" points="105" swimtime="00:03:30.20" resultid="11085" heatid="11728" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.09" />
                    <SPLIT distance="100" swimtime="00:01:34.89" />
                    <SPLIT distance="150" swimtime="00:02:33.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="93" swimtime="00:00:54.99" resultid="11086" heatid="11737" lane="3" entrytime="00:00:56.85" entrycourse="SCM" />
                <RESULT eventid="1331" points="89" swimtime="00:01:49.97" resultid="11087" heatid="11843" lane="6" entrytime="00:01:48.47" entrycourse="SCM" />
                <RESULT eventid="1303" points="106" swimtime="00:01:34.47" resultid="11088" heatid="11824" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Andrade Silva" birthdate="2016-03-15" gender="M" nation="BRA" license="414852" athleteid="11123" externalid="414852">
              <RESULTS>
                <RESULT eventid="1183" points="154" swimtime="00:00:37.58" resultid="11124" heatid="11775" lane="6" entrytime="00:00:41.92" entrycourse="SCM" />
                <RESULT eventid="1137" points="89" swimtime="00:00:48.62" resultid="11125" heatid="11748" lane="2" entrytime="00:01:15.24" entrycourse="SCM" />
                <RESULT eventid="1331" points="126" swimtime="00:01:38.29" resultid="11126" heatid="11843" lane="1" entrytime="00:01:43.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1253" points="124" reactiontime="+89" swimtime="00:00:44.28" resultid="11127" heatid="11802" lane="2" entrytime="00:00:43.55" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elisa" lastname="Damazio Silva" birthdate="2017-01-26" gender="F" nation="BRA" license="421903" athleteid="11146" externalid="421903">
              <RESULTS>
                <RESULT eventid="1324" points="37" swimtime="00:01:08.34" resultid="11147" heatid="11837" lane="4" />
                <RESULT eventid="1258" points="50" swimtime="00:00:32.05" resultid="11148" heatid="11803" lane="3" entrytime="00:00:30.68" entrycourse="SCM" />
                <RESULT eventid="1224" points="30" swimtime="00:00:41.97" resultid="11149" heatid="11785" lane="2" entrytime="00:00:45.24" entrycourse="SCM" />
                <RESULT eventid="1294" points="32" swimtime="00:00:35.05" resultid="11150" heatid="11816" lane="4" entrytime="00:00:37.12" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Debora" lastname="Borges Carneiro" birthdate="1998-05-07" gender="F" nation="BRA" license="266381" athleteid="10895" externalid="266381" level="S14 - SM14">
              <RESULTS>
                <RESULT eventid="1142" points="326" status="EXH" swimtime="00:01:18.51" resultid="10896" heatid="11750" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="527" status="EXH" swimtime="00:01:17.19" resultid="10897" heatid="11791" lane="4" entrytime="00:01:18.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Meneghetti Vidal" birthdate="2015-06-12" gender="M" nation="BRA" license="414851" athleteid="11118" externalid="414851">
              <RESULTS>
                <RESULT eventid="1081" points="133" swimtime="00:03:14.35" resultid="11119" heatid="11729" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.58" />
                    <SPLIT distance="150" swimtime="00:02:27.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1137" points="71" swimtime="00:00:52.48" resultid="11120" heatid="11749" lane="5" entrytime="00:00:48.56" entrycourse="SCM" />
                <RESULT eventid="1331" points="91" reactiontime="+1105" swimtime="00:01:49.18" resultid="11121" heatid="11842" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="133" swimtime="00:01:27.74" resultid="11122" heatid="11825" lane="3" entrytime="00:01:27.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="De Correa" birthdate="2014-12-03" gender="M" nation="BRA" license="403387" athleteid="11069" externalid="403387">
              <RESULTS>
                <RESULT eventid="1152" points="116" swimtime="00:01:37.74" resultid="11070" heatid="11754" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="178" swimtime="00:00:35.83" resultid="11071" heatid="11775" lane="3" entrytime="00:00:36.47" entrycourse="SCM" />
                <RESULT eventid="1303" points="171" swimtime="00:01:20.70" resultid="11072" heatid="11825" lane="4" entrytime="00:01:28.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="160" swimtime="00:03:21.57" resultid="11073" heatid="11847" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.02" />
                    <SPLIT distance="100" swimtime="00:01:38.19" />
                    <SPLIT distance="150" swimtime="00:02:40.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabrielle" lastname="Borba" birthdate="2014-06-15" gender="F" nation="BRA" license="385705" athleteid="10996" externalid="385705">
              <RESULTS>
                <RESULT eventid="1112" points="132" reactiontime="+69" swimtime="00:01:47.55" resultid="10997" heatid="11739" lane="2" />
                <RESULT eventid="1178" points="207" swimtime="00:00:38.73" resultid="10998" heatid="11771" lane="6" entrytime="00:00:40.19" entrycourse="SCM" />
                <RESULT comment="SW 7.2 - Movimentos dos braços não simultâneos.&#10;&#10;&#10;&#10;&#10;&#10;&#10;  (Tempo: 16:38)" eventid="1228" status="DSQ" swimtime="00:01:52.32" resultid="10999" heatid="11789" lane="1" entrytime="00:01:57.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="167" swimtime="00:03:41.22" resultid="11000" heatid="11844" lane="5" entrytime="00:03:58.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.08" />
                    <SPLIT distance="100" swimtime="00:01:51.99" />
                    <SPLIT distance="150" swimtime="00:02:50.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Otavio Luz" birthdate="2013-07-27" gender="M" nation="BRA" license="392111" athleteid="11029" externalid="392111">
              <RESULTS>
                <RESULT eventid="1152" points="173" swimtime="00:01:25.71" resultid="11030" heatid="11755" lane="4" entrytime="00:01:28.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="218" swimtime="00:02:44.93" resultid="11031" heatid="11729" lane="4" entrytime="00:02:53.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                    <SPLIT distance="100" swimtime="00:01:20.47" />
                    <SPLIT distance="150" swimtime="00:02:05.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="210" swimtime="00:01:15.33" resultid="11032" heatid="11826" lane="3" entrytime="00:01:16.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="124" swimtime="00:01:50.58" resultid="11033" heatid="11794" lane="6" entrytime="00:01:55.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Livia" lastname="Rafaela Sita" birthdate="2015-08-10" gender="F" nation="BRA" license="421959" athleteid="11211" externalid="421959">
              <RESULTS>
                <RESULT eventid="1076" points="67" swimtime="00:04:30.84" resultid="11212" heatid="11727" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.61" />
                    <SPLIT distance="150" swimtime="00:03:36.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="152" swimtime="00:00:42.88" resultid="11213" heatid="11770" lane="6" entrytime="00:00:46.61" entrycourse="SCM" />
                <RESULT eventid="1298" points="142" swimtime="00:01:36.25" resultid="11214" heatid="11821" lane="1" entrytime="00:01:45.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="118" reactiontime="+77" swimtime="00:00:51.38" resultid="11215" heatid="11799" lane="3" entrytime="00:00:54.05" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Mochiutti Carneiro" birthdate="2010-04-22" gender="F" nation="BRA" license="370670" athleteid="10942" externalid="370670">
              <RESULTS>
                <RESULT eventid="1060" points="439" swimtime="00:02:25.07" resultid="10943" heatid="11723" lane="2" entrytime="00:02:21.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                    <SPLIT distance="100" swimtime="00:01:09.79" />
                    <SPLIT distance="150" swimtime="00:01:47.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="283" swimtime="00:03:02.10" resultid="10944" heatid="11812" lane="4" entrytime="00:02:54.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                    <SPLIT distance="100" swimtime="00:01:27.43" />
                    <SPLIT distance="150" swimtime="00:02:15.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Tomazeli" birthdate="2017-11-30" gender="M" nation="BRA" license="421901" athleteid="11136" externalid="421901">
              <RESULTS>
                <RESULT eventid="1326" points="55" swimtime="00:00:52.86" resultid="11137" heatid="11840" lane="2" entrytime="00:00:58.84" entrycourse="SCM" />
                <RESULT eventid="1226" points="49" swimtime="00:00:31.23" resultid="11138" heatid="11787" lane="2" />
                <RESULT eventid="1260" points="47" swimtime="00:00:28.53" resultid="11139" heatid="11806" lane="2" entrytime="00:00:31.54" entrycourse="SCM" />
                <RESULT eventid="1296" points="34" swimtime="00:00:30.33" resultid="11140" heatid="11818" lane="2" entrytime="00:00:33.04" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Arthur Da Silva Ortiz" birthdate="2015-04-20" gender="M" nation="BRA" license="399733" athleteid="11059" externalid="399733">
              <RESULTS>
                <RESULT eventid="1081" points="140" swimtime="00:03:11.12" resultid="11060" heatid="11729" lane="2" entrytime="00:03:24.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                    <SPLIT distance="100" swimtime="00:01:32.06" />
                    <SPLIT distance="150" swimtime="00:02:22.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="120" swimtime="00:00:50.51" resultid="11061" heatid="11738" lane="4" entrytime="00:00:48.59" entrycourse="SCM" />
                <RESULT eventid="1331" points="123" swimtime="00:01:38.91" resultid="11062" heatid="11843" lane="4" entrytime="00:01:34.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="151" swimtime="00:01:24.15" resultid="11063" heatid="11826" lane="6" entrytime="00:01:26.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Garcia Cavalcante" birthdate="2011-11-21" gender="M" nation="BRA" license="378200" athleteid="10887" externalid="378200">
              <RESULTS>
                <RESULT eventid="1094" points="359" swimtime="00:02:49.02" resultid="10888" heatid="11732" lane="4" entrytime="00:03:06.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.88" />
                    <SPLIT distance="100" swimtime="00:01:23.67" />
                    <SPLIT distance="150" swimtime="00:02:07.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="350" swimtime="00:01:18.38" resultid="10889" heatid="11796" lane="2" entrytime="00:01:21.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luara" lastname="Polizeli Marostica" birthdate="2017-04-12" gender="F" nation="BRA" license="421958" athleteid="11206" externalid="421958">
              <RESULTS>
                <RESULT eventid="1324" points="19" swimtime="00:01:24.49" resultid="11207" heatid="11838" lane="6" />
                <RESULT eventid="1258" points="47" swimtime="00:00:32.79" resultid="11208" heatid="11803" lane="4" />
                <RESULT eventid="1224" points="34" swimtime="00:00:40.68" resultid="11209" heatid="11785" lane="4" entrytime="00:00:36.95" entrycourse="SCM" />
                <RESULT eventid="1294" points="16" swimtime="00:00:44.27" resultid="11210" heatid="11816" lane="3" entrytime="00:00:36.60" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Corsine Ferreira" birthdate="2010-03-10" gender="F" nation="BRA" license="353591" athleteid="10939" externalid="353591">
              <RESULTS>
                <RESULT eventid="1112" points="326" reactiontime="+75" swimtime="00:01:19.73" resultid="10940" heatid="11742" lane="5" entrytime="00:01:14.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1262" points="326" reactiontime="+69" swimtime="00:02:52.78" resultid="10941" heatid="11808" lane="4" entrytime="00:02:44.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.80" />
                    <SPLIT distance="100" swimtime="00:01:23.69" />
                    <SPLIT distance="150" swimtime="00:02:08.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Forti Francisco" birthdate="2015-07-08" gender="M" nation="BRA" license="392104" athleteid="11011" externalid="392104">
              <RESULTS>
                <RESULT eventid="1081" points="112" swimtime="00:03:25.76" resultid="11012" heatid="11728" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.12" />
                    <SPLIT distance="100" swimtime="00:01:30.21" />
                    <SPLIT distance="150" swimtime="00:02:29.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="97" swimtime="00:00:54.23" resultid="11013" heatid="11738" lane="6" entrytime="00:00:56.39" entrycourse="SCM" />
                <RESULT eventid="1331" points="104" swimtime="00:01:44.69" resultid="11014" heatid="11842" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="103" swimtime="00:01:35.54" resultid="11015" heatid="11825" lane="2" entrytime="00:01:33.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Pacheco" birthdate="2006-12-20" gender="M" nation="BRA" license="336850" athleteid="10901" externalid="336850">
              <RESULTS>
                <RESULT eventid="1152" points="453" swimtime="00:01:02.17" resultid="10902" heatid="11758" lane="1" entrytime="00:01:02.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="414" swimtime="00:02:23.33" resultid="10903" heatid="11815" lane="2" entrytime="00:02:21.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                    <SPLIT distance="100" swimtime="00:01:06.86" />
                    <SPLIT distance="150" swimtime="00:01:44.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Eduardo Ebiner" birthdate="2013-07-29" gender="M" nation="BRA" license="397371" athleteid="11054" externalid="397371">
              <RESULTS>
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Tempo: 11:21), Na volta dos 25m." eventid="1152" status="DSQ" swimtime="00:01:47.21" resultid="11055" heatid="11754" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="160" swimtime="00:00:37.10" resultid="11056" heatid="11775" lane="2" entrytime="00:00:37.85" entrycourse="SCM" />
                <RESULT eventid="1238" points="137" swimtime="00:01:47.20" resultid="11057" heatid="11793" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1214" points="157" swimtime="00:06:32.70" resultid="11058" heatid="11781" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.76" />
                    <SPLIT distance="100" swimtime="00:01:33.13" />
                    <SPLIT distance="150" swimtime="00:02:22.89" />
                    <SPLIT distance="200" swimtime="00:03:11.67" />
                    <SPLIT distance="250" swimtime="00:04:00.71" />
                    <SPLIT distance="300" swimtime="00:04:51.41" />
                    <SPLIT distance="350" swimtime="00:05:42.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietro" lastname="Nabas De Assis" birthdate="2011-07-09" gender="M" nation="BRA" license="366968" athleteid="10932" externalid="366968">
              <RESULTS>
                <RESULT comment="SW 5.3 - Totalmente submerso durante o nado." eventid="1170" status="DSQ" swimtime="00:00:36.93" resultid="10933" heatid="11765" lane="3" entrytime="00:00:29.68" entrycourse="SCM" />
                <RESULT eventid="1238" points="386" swimtime="00:01:15.87" resultid="10934" heatid="11797" lane="6" entrytime="00:01:16.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnes" lastname="Sophie Amadei" birthdate="2014-01-10" gender="F" nation="BRA" license="403388" athleteid="11074" externalid="403388">
              <RESULTS>
                <RESULT eventid="1142" points="104" swimtime="00:01:54.91" resultid="11075" heatid="11750" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="195" swimtime="00:00:39.48" resultid="11076" heatid="11771" lane="1" entrytime="00:00:39.86" entrycourse="SCM" />
                <RESULT eventid="1204" points="152" swimtime="00:07:13.12" resultid="11077" heatid="11779" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.53" />
                    <SPLIT distance="100" swimtime="00:01:40.94" />
                    <SPLIT distance="150" swimtime="00:02:38.22" />
                    <SPLIT distance="200" swimtime="00:03:32.79" />
                    <SPLIT distance="250" swimtime="00:04:28.96" />
                    <SPLIT distance="300" swimtime="00:05:26.32" />
                    <SPLIT distance="350" swimtime="00:06:20.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="127" reactiontime="+48" swimtime="00:00:50.16" resultid="11078" heatid="11799" lane="4" entrytime="00:00:56.96" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wellington" lastname="De Lima" birthdate="2008-03-01" gender="M" nation="BRA" license="370024" athleteid="10876" externalid="370024">
              <RESULTS>
                <RESULT eventid="1122" points="392" swimtime="00:01:06.02" resultid="10877" heatid="11746" lane="4" entrytime="00:01:07.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1316" points="530" swimtime="00:00:55.39" resultid="10878" heatid="11836" lane="2" entrytime="00:00:55.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1214" points="454" swimtime="00:04:36.05" resultid="10879" heatid="11781" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.46" />
                    <SPLIT distance="100" swimtime="00:01:01.95" />
                    <SPLIT distance="150" swimtime="00:01:36.31" />
                    <SPLIT distance="200" swimtime="00:02:11.59" />
                    <SPLIT distance="250" swimtime="00:02:47.75" />
                    <SPLIT distance="300" swimtime="00:03:23.78" />
                    <SPLIT distance="350" swimtime="00:03:59.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15981" nation="BRA" region="PR" clubid="10839" name="Quinto Nado" shortname="5º Nado">
          <ATHLETES>
            <ATHLETE firstname="Laura" lastname="Takemura Couto" birthdate="2010-02-08" gender="F" nation="BRA" license="376950" athleteid="10850" externalid="376950">
              <RESULTS>
                <RESULT eventid="1142" points="456" swimtime="00:01:10.20" resultid="10851" heatid="11752" lane="6" entrytime="00:01:22.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="554" swimtime="00:02:14.30" resultid="10852" heatid="11723" lane="4" entrytime="00:02:13.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                    <SPLIT distance="100" swimtime="00:01:05.52" />
                    <SPLIT distance="150" swimtime="00:01:40.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1308" points="530" swimtime="00:01:02.06" resultid="10853" heatid="11830" lane="3" entrytime="00:01:00.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1262" points="412" reactiontime="+67" swimtime="00:02:39.72" resultid="10854" heatid="11808" lane="5" entrytime="00:02:50.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                    <SPLIT distance="100" swimtime="00:01:18.87" />
                    <SPLIT distance="150" swimtime="00:01:59.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Poletti Veiga" birthdate="2010-10-01" gender="F" nation="BRA" license="376951" athleteid="10845" externalid="376951">
              <RESULTS>
                <RESULT eventid="1060" points="560" swimtime="00:02:13.79" resultid="10846" heatid="11723" lane="3" entrytime="00:02:12.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                    <SPLIT distance="100" swimtime="00:01:05.39" />
                    <SPLIT distance="150" swimtime="00:01:39.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="491" swimtime="00:10:04.84" resultid="10847" heatid="11777" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:13.65" />
                    <SPLIT distance="150" swimtime="00:01:52.62" />
                    <SPLIT distance="200" swimtime="00:02:31.53" />
                    <SPLIT distance="250" swimtime="00:03:10.90" />
                    <SPLIT distance="300" swimtime="00:03:49.73" />
                    <SPLIT distance="350" swimtime="00:04:29.02" />
                    <SPLIT distance="400" swimtime="00:05:07.06" />
                    <SPLIT distance="450" swimtime="00:05:45.38" />
                    <SPLIT distance="500" swimtime="00:06:23.57" />
                    <SPLIT distance="550" swimtime="00:07:01.44" />
                    <SPLIT distance="600" swimtime="00:07:38.78" />
                    <SPLIT distance="650" swimtime="00:08:16.06" />
                    <SPLIT distance="700" swimtime="00:08:53.26" />
                    <SPLIT distance="750" swimtime="00:09:29.60" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.1 - Mais de uma pernada de borboleta antes da primeira pernada de peito após o início ou a virada.  (Tempo: 19:36), Após a volta dos 100m (Peito, Medley Individual)." eventid="1334" status="DSQ" swimtime="00:02:45.28" resultid="10848" heatid="11845" lane="4" entrytime="00:02:48.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                    <SPLIT distance="100" swimtime="00:01:18.82" />
                    <SPLIT distance="150" swimtime="00:02:10.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="488" swimtime="00:04:53.62" resultid="10849" heatid="11780" lane="3" entrytime="00:04:45.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                    <SPLIT distance="100" swimtime="00:01:09.81" />
                    <SPLIT distance="150" swimtime="00:01:47.13" />
                    <SPLIT distance="200" swimtime="00:02:24.38" />
                    <SPLIT distance="250" swimtime="00:03:01.61" />
                    <SPLIT distance="300" swimtime="00:03:39.26" />
                    <SPLIT distance="350" swimtime="00:04:16.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Kikuchi Fujii" birthdate="2007-01-04" gender="M" nation="BRA" license="297805" athleteid="10840" externalid="297805">
              <RESULTS>
                <RESULT eventid="1152" points="576" swimtime="00:00:57.40" resultid="10841" heatid="11754" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1094" points="600" swimtime="00:02:22.43" resultid="10842" heatid="11733" lane="3" entrytime="00:02:19.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                    <SPLIT distance="100" swimtime="00:01:08.98" />
                    <SPLIT distance="150" swimtime="00:01:45.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="601" swimtime="00:01:05.49" resultid="10843" heatid="11797" lane="3" entrytime="00:01:03.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="458" swimtime="00:02:18.55" resultid="10844" heatid="11814" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                    <SPLIT distance="100" swimtime="00:01:05.76" />
                    <SPLIT distance="150" swimtime="00:01:42.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco" lastname="Silva Telles" birthdate="2011-07-19" gender="M" nation="BRA" license="377311" athleteid="10855" externalid="377311">
              <RESULTS>
                <RESULT eventid="1094" points="296" swimtime="00:03:00.13" resultid="10856" heatid="11732" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.97" />
                    <SPLIT distance="100" swimtime="00:01:26.68" />
                    <SPLIT distance="150" swimtime="00:02:15.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="289" swimtime="00:00:30.47" resultid="10857" heatid="11765" lane="6" entrytime="00:00:32.28" entrycourse="SCM" />
                <RESULT eventid="1316" points="298" swimtime="00:01:07.11" resultid="10858" heatid="11831" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente., Na volta dos 75m." eventid="1238" status="DSQ" swimtime="00:01:20.76" resultid="10859" heatid="11796" lane="1" entrytime="00:01:24.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Fernanda Iossaqui" birthdate="2014-08-01" gender="F" nation="BRA" license="421517" athleteid="10860" externalid="421517">
              <RESULTS>
                <RESULT eventid="1178" points="173" swimtime="00:00:41.11" resultid="10861" heatid="11770" lane="3" entrytime="00:00:41.65" entrycourse="SCM" />
                <RESULT eventid="1102" points="145" swimtime="00:00:53.98" resultid="10862" heatid="11734" lane="2" />
                <RESULT eventid="1298" points="161" swimtime="00:01:32.26" resultid="10863" heatid="11819" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="156" swimtime="00:01:55.82" resultid="10864" heatid="11788" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15969" nation="BRA" region="RJ" clubid="11381" name="Estados Unidos Da América" shortname="Eua">
          <ATHLETES>
            <ATHLETE firstname="Sophia" lastname="Alanis Whitney" birthdate="2007-07-21" gender="F" nation="USA" license="V397028" athleteid="11382" externalid="V397028">
              <RESULTS>
                <RESULT eventid="1142" points="518" status="EXH" swimtime="00:01:07.30" resultid="11383" heatid="11752" lane="3" entrytime="00:01:05.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="477" reactiontime="+75" status="EXH" swimtime="00:01:10.24" resultid="11384" heatid="11742" lane="3" entrytime="00:01:11.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="448" status="EXH" swimtime="00:02:36.28" resultid="11385" heatid="11812" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                    <SPLIT distance="100" swimtime="00:01:13.16" />
                    <SPLIT distance="150" swimtime="00:01:53.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="434" status="EXH" swimtime="00:02:40.83" resultid="11386" heatid="11844" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                    <SPLIT distance="100" swimtime="00:01:15.10" />
                    <SPLIT distance="150" swimtime="00:02:05.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16053" nation="BRA" region="PR" clubid="11387" name="Fábrica De Nadadores" shortname="Fábrica">
          <ATHLETES>
            <ATHLETE firstname="Victor" lastname="Kenji Yamaguchi" birthdate="2011-08-25" gender="M" nation="BRA" license="385708" athleteid="11431" externalid="385708">
              <RESULTS>
                <RESULT eventid="1152" points="333" swimtime="00:01:08.93" resultid="11432" heatid="11756" lane="2" entrytime="00:01:12.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="322" swimtime="00:02:35.85" resultid="11433" heatid="11813" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                    <SPLIT distance="100" swimtime="00:01:14.22" />
                    <SPLIT distance="150" swimtime="00:01:55.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="309" swimtime="00:02:42.06" resultid="11434" heatid="11849" lane="2" entrytime="00:02:41.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                    <SPLIT distance="100" swimtime="00:01:17.31" />
                    <SPLIT distance="150" swimtime="00:02:05.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Ognibeni Paupitz" birthdate="2014-08-08" gender="F" nation="BRA" license="406923" athleteid="11518" externalid="406923">
              <RESULTS>
                <RESULT eventid="1178" points="190" swimtime="00:00:39.88" resultid="11519" heatid="11770" lane="2" entrytime="00:00:43.36" entrycourse="SCM" />
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Tempo: 10:19), Na volta dos 25m." eventid="1102" status="DSQ" swimtime="00:00:51.80" resultid="11520" heatid="11736" lane="5" entrytime="00:00:55.61" entrycourse="SCM" />
                <RESULT eventid="1298" points="136" swimtime="00:01:37.69" resultid="11521" heatid="11821" lane="6" entrytime="00:01:54.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="144" swimtime="00:01:58.79" resultid="11522" heatid="11788" lane="3" entrytime="00:02:09.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Tiemi Yamaguchi" birthdate="2013-02-28" gender="F" nation="BRA" license="385707" athleteid="11467" externalid="385707">
              <RESULTS>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Tempo: 11:08)" eventid="1142" status="DSQ" swimtime="00:01:20.91" resultid="11468" heatid="11751" lane="2" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.62" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 6.4 - A virada não foi iniciada após a conclusão do movimento de braço, após sair da posição de costas.  (Tempo: 10:30), Na volta dos 50m." eventid="1112" reactiontime="+67" status="DSQ" swimtime="00:01:20.96" resultid="11469" heatid="11739" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="300" swimtime="00:01:15.04" resultid="11470" heatid="11822" lane="2" entrytime="00:01:17.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="331" swimtime="00:05:34.21" resultid="11471" heatid="11780" lane="1" entrytime="00:05:42.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                    <SPLIT distance="100" swimtime="00:01:17.64" />
                    <SPLIT distance="150" swimtime="00:02:00.79" />
                    <SPLIT distance="200" swimtime="00:02:44.12" />
                    <SPLIT distance="250" swimtime="00:03:27.60" />
                    <SPLIT distance="300" swimtime="00:04:10.62" />
                    <SPLIT distance="350" swimtime="00:04:52.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Miranda Amorim" birthdate="2016-02-06" gender="F" nation="BRA" license="421991" athleteid="11550" externalid="421991">
              <RESULTS>
                <RESULT eventid="1178" points="85" swimtime="00:00:52.01" resultid="11551" heatid="11768" lane="4" entrytime="00:00:57.91" entrycourse="SCM" />
                <RESULT eventid="1102" points="94" swimtime="00:01:02.32" resultid="11552" heatid="11735" lane="2" entrytime="00:01:05.90" entrycourse="SCM" />
                <RESULT eventid="1298" status="DNS" swimtime="00:00:00.00" resultid="11553" heatid="11820" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Jupi Takaki" birthdate="2013-03-26" gender="F" nation="BRA" license="391845" athleteid="11477" externalid="391845">
              <RESULTS>
                <RESULT eventid="1142" points="282" swimtime="00:01:22.33" resultid="11478" heatid="11751" lane="1" entrytime="00:01:27.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1076" points="330" swimtime="00:02:39.53" resultid="11479" heatid="11727" lane="3" entrytime="00:02:46.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                    <SPLIT distance="100" swimtime="00:01:17.78" />
                    <SPLIT distance="150" swimtime="00:01:59.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="307" swimtime="00:01:14.47" resultid="11480" heatid="11821" lane="3" entrytime="00:01:20.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="300" swimtime="00:05:45.24" resultid="11481" heatid="11780" lane="6" entrytime="00:05:56.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.43" />
                    <SPLIT distance="100" swimtime="00:01:20.05" />
                    <SPLIT distance="150" swimtime="00:02:04.28" />
                    <SPLIT distance="200" swimtime="00:02:48.98" />
                    <SPLIT distance="250" swimtime="00:03:34.23" />
                    <SPLIT distance="300" swimtime="00:04:18.44" />
                    <SPLIT distance="350" swimtime="00:05:02.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kauana" lastname="De Leal" birthdate="2016-02-20" gender="F" nation="BRA" license="417997" athleteid="11541" externalid="417997">
              <RESULTS>
                <RESULT eventid="1178" points="39" swimtime="00:01:07.16" resultid="11542" heatid="11768" lane="1" entrytime="00:01:11.44" entrycourse="SCM" />
                <RESULT eventid="1102" points="57" swimtime="00:01:13.59" resultid="11543" heatid="11734" lane="4" entrytime="00:01:30.54" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Livia" lastname="Eloisa Silva" birthdate="2012-03-03" gender="F" nation="BRA" license="399725" athleteid="11505" externalid="399725">
              <RESULTS>
                <RESULT eventid="1060" points="163" swimtime="00:03:21.57" resultid="11506" heatid="11722" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.27" />
                    <SPLIT distance="100" swimtime="00:01:36.01" />
                    <SPLIT distance="150" swimtime="00:02:28.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1162" points="170" swimtime="00:00:41.39" resultid="11507" heatid="11759" lane="2" entrytime="00:00:47.16" entrycourse="SCM" />
                <RESULT eventid="1308" points="183" swimtime="00:01:28.38" resultid="11508" heatid="11827" lane="3" entrytime="00:01:43.89" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Dias Rezende" birthdate="2016-03-04" gender="F" nation="BRA" license="406929" athleteid="11530" externalid="406929">
              <RESULTS>
                <RESULT eventid="1178" status="DNS" swimtime="00:00:00.00" resultid="11531" heatid="11768" lane="5" entrytime="00:01:08.48" entrycourse="SCM" />
                <RESULT eventid="1102" status="DNS" swimtime="00:00:00.00" resultid="11532" heatid="11734" lane="3" entrytime="00:01:19.05" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eloah" lastname="Juvedi Trindade" birthdate="2011-03-05" gender="F" nation="BRA" license="396829" athleteid="11492" externalid="396829">
              <RESULTS>
                <RESULT eventid="1142" points="212" swimtime="00:01:30.56" resultid="11493" heatid="11750" lane="3" entrytime="00:01:42.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1162" points="343" swimtime="00:00:32.73" resultid="11494" heatid="11760" lane="5" entrytime="00:00:33.38" entrycourse="SCM" />
                <RESULT eventid="1308" points="329" swimtime="00:01:12.78" resultid="11495" heatid="11828" lane="3" entrytime="00:01:16.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="266" swimtime="00:03:09.28" resultid="11496" heatid="11844" lane="4" entrytime="00:03:29.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.89" />
                    <SPLIT distance="100" swimtime="00:01:33.63" />
                    <SPLIT distance="150" swimtime="00:02:28.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eloah" lastname="Frasson" birthdate="2012-06-14" gender="F" nation="BRA" license="378338" athleteid="11447" externalid="378338">
              <RESULTS>
                <RESULT eventid="1086" points="307" swimtime="00:03:19.45" resultid="11448" heatid="11731" lane="6" entrytime="00:03:20.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.45" />
                    <SPLIT distance="100" swimtime="00:01:33.67" />
                    <SPLIT distance="150" swimtime="00:02:26.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1162" points="339" swimtime="00:00:32.88" resultid="11449" heatid="11760" lane="6" entrytime="00:00:35.49" entrycourse="SCM" />
                <RESULT eventid="1308" points="338" swimtime="00:01:12.10" resultid="11450" heatid="11828" lane="2" entrytime="00:01:18.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="375" swimtime="00:01:26.40" resultid="11451" heatid="11790" lane="2" entrytime="00:01:27.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marco" lastname="Manzotti Marchi" birthdate="2015-06-26" gender="M" nation="BRA" license="396849" athleteid="11497" externalid="396849">
              <RESULTS>
                <RESULT eventid="1137" status="DNS" swimtime="00:00:00.00" resultid="11498" heatid="11749" lane="2" entrytime="00:00:46.57" entrycourse="SCM" />
                <RESULT eventid="1331" status="DNS" swimtime="00:00:00.00" resultid="11499" heatid="11842" lane="1" />
                <RESULT eventid="1303" status="DNS" swimtime="00:00:00.00" resultid="11500" heatid="11825" lane="1" entrytime="00:01:35.45" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Donatello" lastname="Dacome" birthdate="2015-08-24" gender="M" nation="BRA" license="421988" athleteid="11547" externalid="421988">
              <RESULTS>
                <RESULT eventid="1183" points="29" swimtime="00:01:05.55" resultid="11548" heatid="11773" lane="5" />
                <RESULT eventid="1107" points="57" swimtime="00:01:04.48" resultid="11549" heatid="11737" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="Jacobsen Donati" birthdate="2011-07-14" gender="M" nation="BRA" license="391851" athleteid="11426" externalid="391851">
              <RESULTS>
                <RESULT eventid="1152" points="377" swimtime="00:01:06.09" resultid="11427" heatid="11757" lane="6" entrytime="00:01:09.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="454" swimtime="00:02:09.28" resultid="11428" heatid="11725" lane="1" entrytime="00:02:17.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.41" />
                    <SPLIT distance="100" swimtime="00:01:01.56" />
                    <SPLIT distance="150" swimtime="00:01:35.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="394" swimtime="00:02:29.51" resultid="11429" heatid="11846" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                    <SPLIT distance="100" swimtime="00:01:07.81" />
                    <SPLIT distance="150" swimtime="00:01:56.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1214" points="401" swimtime="00:04:47.68" resultid="11430" heatid="11783" lane="5" entrytime="00:04:57.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.91" />
                    <SPLIT distance="100" swimtime="00:01:06.91" />
                    <SPLIT distance="150" swimtime="00:01:42.89" />
                    <SPLIT distance="200" swimtime="00:02:19.64" />
                    <SPLIT distance="250" swimtime="00:02:56.49" />
                    <SPLIT distance="300" swimtime="00:03:33.69" />
                    <SPLIT distance="350" swimtime="00:04:10.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theodoro" lastname="Marques Serra" birthdate="2009-11-24" gender="M" nation="BRA" license="370661" athleteid="11411" externalid="370661">
              <RESULTS>
                <RESULT eventid="1068" points="471" swimtime="00:02:07.68" resultid="11412" heatid="11726" lane="6" entrytime="00:02:10.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                    <SPLIT distance="100" swimtime="00:01:01.33" />
                    <SPLIT distance="150" swimtime="00:01:35.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="425" swimtime="00:09:45.69" resultid="11413" heatid="11778" lane="3" entrytime="00:10:18.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                    <SPLIT distance="100" swimtime="00:01:08.10" />
                    <SPLIT distance="150" swimtime="00:01:45.60" />
                    <SPLIT distance="200" swimtime="00:02:23.24" />
                    <SPLIT distance="250" swimtime="00:03:01.10" />
                    <SPLIT distance="300" swimtime="00:03:38.09" />
                    <SPLIT distance="350" swimtime="00:04:15.85" />
                    <SPLIT distance="400" swimtime="00:04:53.84" />
                    <SPLIT distance="450" swimtime="00:05:31.15" />
                    <SPLIT distance="500" swimtime="00:06:08.63" />
                    <SPLIT distance="550" swimtime="00:06:44.96" />
                    <SPLIT distance="600" swimtime="00:07:21.33" />
                    <SPLIT distance="650" swimtime="00:07:58.39" />
                    <SPLIT distance="700" swimtime="00:08:35.06" />
                    <SPLIT distance="750" swimtime="00:09:11.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="253" swimtime="00:02:48.90" resultid="11414" heatid="11813" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                    <SPLIT distance="100" swimtime="00:01:17.79" />
                    <SPLIT distance="150" swimtime="00:02:03.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1214" points="437" swimtime="00:04:39.55" resultid="11415" heatid="11783" lane="2" entrytime="00:04:37.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                    <SPLIT distance="100" swimtime="00:01:03.78" />
                    <SPLIT distance="150" swimtime="00:01:39.36" />
                    <SPLIT distance="200" swimtime="00:02:15.74" />
                    <SPLIT distance="250" swimtime="00:02:52.03" />
                    <SPLIT distance="300" swimtime="00:03:28.24" />
                    <SPLIT distance="350" swimtime="00:04:04.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Silveira De Almeida" birthdate="2008-07-08" gender="M" nation="BRA" license="368152" athleteid="11440" externalid="368152">
              <RESULTS>
                <RESULT eventid="1152" points="373" swimtime="00:01:06.34" resultid="11441" heatid="11758" lane="5" entrytime="00:01:01.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="344" swimtime="00:02:21.76" resultid="11442" heatid="11724" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                    <SPLIT distance="100" swimtime="00:01:05.06" />
                    <SPLIT distance="150" swimtime="00:01:43.27" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 5.3 - Totalmente submerso durante o nado.  (Tempo: 18:48)" eventid="1316" status="DSQ" swimtime="00:01:10.31" resultid="11443" heatid="11831" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="345" swimtime="00:02:32.33" resultid="11444" heatid="11815" lane="4" entrytime="00:02:17.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:01:51.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Moreschi" birthdate="2012-08-09" gender="M" nation="BRA" license="385715" athleteid="11421" externalid="385715">
              <RESULTS>
                <RESULT eventid="1152" points="176" swimtime="00:01:25.23" resultid="11422" heatid="11755" lane="3" entrytime="00:01:25.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1094" points="256" swimtime="00:03:09.08" resultid="11423" heatid="11732" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                    <SPLIT distance="100" swimtime="00:01:31.86" />
                    <SPLIT distance="150" swimtime="00:02:21.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="242" swimtime="00:01:28.61" resultid="11424" heatid="11794" lane="3" entrytime="00:01:35.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="178" swimtime="00:03:09.93" resultid="11425" heatid="11814" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.53" />
                    <SPLIT distance="100" swimtime="00:01:30.29" />
                    <SPLIT distance="150" swimtime="00:02:21.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Schmeiske Ruivo" birthdate="2013-10-21" gender="F" nation="BRA" license="402006" athleteid="11509" externalid="402006">
              <RESULTS>
                <RESULT eventid="1132" points="295" swimtime="00:00:36.62" resultid="11510" heatid="11747" lane="3" entrytime="00:00:35.01" entrycourse="SCM" />
                <RESULT eventid="1178" points="436" swimtime="00:00:30.22" resultid="11511" heatid="11772" lane="4" entrytime="00:00:30.68" entrycourse="SCM" />
                <RESULT eventid="1298" points="384" swimtime="00:01:09.08" resultid="11512" heatid="11822" lane="1" entrytime="00:01:19.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="383" swimtime="00:01:25.86" resultid="11513" heatid="11790" lane="6" entrytime="00:01:30.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Britto" birthdate="2012-10-04" gender="M" nation="BRA" license="378350" athleteid="11402" externalid="378350">
              <RESULTS>
                <RESULT eventid="1152" points="215" swimtime="00:01:19.65" resultid="11403" heatid="11756" lane="6" entrytime="00:01:25.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1122" points="291" swimtime="00:01:12.85" resultid="11404" heatid="11745" lane="2" entrytime="00:01:18.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="309" reactiontime="+66" swimtime="00:02:36.20" resultid="11405" heatid="11809" lane="4" entrytime="00:02:53.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.31" />
                    <SPLIT distance="100" swimtime="00:01:15.16" />
                    <SPLIT distance="150" swimtime="00:01:56.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elen" lastname="Torres Gomes" birthdate="2015-10-15" gender="F" nation="BRA" license="396850" athleteid="11501" externalid="396850">
              <RESULTS>
                <RESULT eventid="1102" points="104" swimtime="00:01:00.20" resultid="11502" heatid="11735" lane="4" entrytime="00:01:03.23" entrycourse="SCM" />
                <RESULT eventid="1328" points="99" swimtime="00:02:01.86" resultid="11503" heatid="11841" lane="3" entrytime="00:02:04.07" entrycourse="SCM" />
                <RESULT eventid="1298" points="107" swimtime="00:01:45.57" resultid="11504" heatid="11821" lane="5" entrytime="00:01:41.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dante" lastname="Gabriel Rossi" birthdate="2016-01-19" gender="M" nation="BRA" license="406928" athleteid="11526" externalid="406928">
              <RESULTS>
                <RESULT eventid="1183" points="102" swimtime="00:00:43.12" resultid="11527" heatid="11774" lane="3" entrytime="00:00:44.61" entrycourse="SCM" />
                <RESULT eventid="1137" points="71" swimtime="00:00:52.45" resultid="11528" heatid="11748" lane="4" entrytime="00:01:03.18" entrycourse="SCM" />
                <RESULT eventid="1253" points="75" reactiontime="+60" swimtime="00:00:52.28" resultid="11529" heatid="11801" lane="2" entrytime="00:00:54.19" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Bagatim" birthdate="2014-05-27" gender="F" nation="BRA" license="378353" athleteid="11457" externalid="378353">
              <RESULTS>
                <RESULT eventid="1132" points="322" swimtime="00:00:35.56" resultid="11458" heatid="11747" lane="4" entrytime="00:00:35.89" entrycourse="SCM" />
                <RESULT eventid="1178" points="300" swimtime="00:00:34.22" resultid="11459" heatid="11772" lane="5" entrytime="00:00:34.23" entrycourse="SCM" />
                <RESULT eventid="1298" points="293" swimtime="00:01:15.59" resultid="11460" heatid="11822" lane="6" entrytime="00:01:19.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="227" swimtime="00:01:42.20" resultid="11461" heatid="11788" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Harada Otero" birthdate="2014-11-06" gender="M" nation="BRA" license="424615" athleteid="11565" externalid="424615">
              <RESULTS>
                <RESULT eventid="1122" points="72" reactiontime="+131" swimtime="00:01:55.78" resultid="11566" heatid="11743" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="72" swimtime="00:00:48.37" resultid="11567" heatid="11773" lane="2" />
                <RESULT eventid="1303" points="62" swimtime="00:01:52.85" resultid="11568" heatid="11824" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1253" points="59" reactiontime="+124" swimtime="00:00:56.51" resultid="11569" heatid="11801" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruna" lastname="Mine Moreschi" birthdate="2017-11-15" gender="F" nation="BRA" license="421987" athleteid="11544" externalid="421987">
              <RESULTS>
                <RESULT eventid="1324" points="27" swimtime="00:01:15.67" resultid="11545" heatid="11837" lane="2" />
                <RESULT eventid="1224" points="30" swimtime="00:00:41.99" resultid="11546" heatid="11784" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Valentina Gozaga" birthdate="2014-06-28" gender="F" nation="BRA" license="385709" athleteid="11472" externalid="385709">
              <RESULTS>
                <RESULT eventid="1178" points="237" swimtime="00:00:37.01" resultid="11473" heatid="11771" lane="5" entrytime="00:00:39.26" entrycourse="SCM" />
                <RESULT eventid="1102" points="186" swimtime="00:00:49.65" resultid="11474" heatid="11736" lane="4" entrytime="00:00:53.53" entrycourse="SCM" />
                <RESULT eventid="1228" points="168" swimtime="00:01:53.01" resultid="11475" heatid="11789" lane="6" entrytime="00:01:58.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="163" reactiontime="+72" swimtime="00:00:46.20" resultid="11476" heatid="11800" lane="1" entrytime="00:00:47.44" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Gabriel Iusten" birthdate="2011-04-11" gender="M" nation="BRA" license="406920" athleteid="11514" externalid="406920">
              <RESULTS>
                <RESULT eventid="1170" points="127" swimtime="00:00:40.08" resultid="11515" heatid="11762" lane="4" entrytime="00:00:43.68" entrycourse="SCM" />
                <RESULT eventid="1316" points="121" swimtime="00:01:30.42" resultid="11516" heatid="11831" lane="4" entrytime="00:01:34.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="107" swimtime="00:01:56.23" resultid="11517" heatid="11793" lane="5" entrytime="00:02:09.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Sales" birthdate="2011-02-28" gender="F" nation="BRA" license="374103" athleteid="11445" externalid="374103">
              <RESULTS>
                <RESULT comment="SW 8.5 - Mais de um movimento de braço sob (em baixo) a água após o início ou a virada.&#10;&#10;&#10;&#10;&#10;&#10;&#10;  (Tempo: 19:08)" eventid="1278" status="DSQ" swimtime="00:02:54.35" resultid="11446" heatid="11871" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                    <SPLIT distance="100" swimtime="00:01:16.81" />
                    <SPLIT distance="150" swimtime="00:02:01.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruna" lastname="Scalise Drapzichinski" birthdate="2012-03-07" gender="F" nation="BRA" license="378349" athleteid="11393" externalid="378349">
              <RESULTS>
                <RESULT eventid="1086" points="446" swimtime="00:02:56.09" resultid="11394" heatid="11731" lane="5" entrytime="00:03:06.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.29" />
                    <SPLIT distance="100" swimtime="00:01:22.37" />
                    <SPLIT distance="150" swimtime="00:02:09.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1162" points="444" swimtime="00:00:30.04" resultid="11395" heatid="11761" lane="3" entrytime="00:00:28.70" entrycourse="SCM" />
                <RESULT eventid="1308" points="451" swimtime="00:01:05.49" resultid="11396" heatid="11830" lane="2" entrytime="00:01:07.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="511" swimtime="00:01:17.97" resultid="11397" heatid="11791" lane="3" entrytime="00:01:18.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Limonta Moreto" birthdate="2015-06-29" gender="M" nation="BRA" license="408979" athleteid="11537" externalid="408979">
              <RESULTS>
                <RESULT eventid="1183" points="93" swimtime="00:00:44.39" resultid="11538" heatid="11773" lane="4" />
                <RESULT eventid="1107" points="80" swimtime="00:00:57.75" resultid="11539" heatid="11737" lane="5" />
                <RESULT eventid="1303" points="81" swimtime="00:01:43.48" resultid="11540" heatid="11823" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Rossi" birthdate="2012-05-21" gender="M" nation="BRA" license="378346" athleteid="11452" externalid="378346">
              <RESULTS>
                <RESULT eventid="1122" points="192" swimtime="00:01:23.72" resultid="11453" heatid="11745" lane="6" entrytime="00:01:23.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="319" swimtime="00:00:29.48" resultid="11454" heatid="11765" lane="2" entrytime="00:00:31.19" entrycourse="SCM" />
                <RESULT eventid="1316" points="283" swimtime="00:01:08.22" resultid="11455" heatid="11834" lane="5" entrytime="00:01:10.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="223" swimtime="00:03:00.70" resultid="11456" heatid="11847" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.07" />
                    <SPLIT distance="100" swimtime="00:01:28.39" />
                    <SPLIT distance="150" swimtime="00:02:22.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Traci Rodrigues" birthdate="2014-10-27" gender="M" nation="BRA" license="406926" athleteid="11523" externalid="406926">
              <RESULTS>
                <RESULT eventid="1303" points="120" swimtime="00:01:30.78" resultid="11524" heatid="11825" lane="5" entrytime="00:01:34.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="104" swimtime="00:01:57.34" resultid="11525" heatid="11793" lane="4" entrytime="00:02:04.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Gevaerd Verssutti Garcia" birthdate="2013-10-15" gender="F" nation="BRA" license="378404" athleteid="11462" externalid="378404">
              <RESULTS>
                <RESULT eventid="1142" points="191" swimtime="00:01:33.83" resultid="11463" heatid="11750" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="286" reactiontime="+76" swimtime="00:01:23.31" resultid="11464" heatid="11740" lane="3" entrytime="00:01:27.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="298" swimtime="00:01:15.19" resultid="11465" heatid="11822" lane="5" entrytime="00:01:18.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="260" swimtime="00:06:02.21" resultid="11466" heatid="11779" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.09" />
                    <SPLIT distance="100" swimtime="00:01:24.09" />
                    <SPLIT distance="150" swimtime="00:02:10.53" />
                    <SPLIT distance="200" swimtime="00:02:58.17" />
                    <SPLIT distance="250" swimtime="00:03:45.20" />
                    <SPLIT distance="300" swimtime="00:04:32.29" />
                    <SPLIT distance="350" swimtime="00:05:18.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Ricardo Loureiro" birthdate="2012-07-25" gender="M" nation="BRA" license="424616" athleteid="11570" externalid="424616">
              <RESULTS>
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Tempo: 11:21), Na volta dos 25m, 50m, 75m." eventid="1152" status="DSQ" swimtime="00:01:46.28" resultid="11571" heatid="11754" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="144" swimtime="00:00:38.45" resultid="11572" heatid="11762" lane="2" />
                <RESULT eventid="1316" points="134" swimtime="00:01:27.62" resultid="11573" heatid="11831" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Imai" birthdate="2017-06-28" gender="M" nation="BRA" license="424614" athleteid="11562" externalid="424614">
              <RESULTS>
                <RESULT eventid="1326" points="79" swimtime="00:00:46.90" resultid="11563" heatid="11839" lane="2" />
                <RESULT eventid="1226" points="53" swimtime="00:00:30.37" resultid="11564" heatid="11786" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Braga" birthdate="2010-05-07" gender="M" nation="BRA" license="378345" athleteid="11388" externalid="378345">
              <RESULTS>
                <RESULT eventid="1094" points="480" swimtime="00:02:33.39" resultid="11389" heatid="11733" lane="4" entrytime="00:02:37.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.20" />
                    <SPLIT distance="100" swimtime="00:01:15.03" />
                    <SPLIT distance="150" swimtime="00:01:55.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="321" swimtime="00:10:42.87" resultid="11390" heatid="11778" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                    <SPLIT distance="100" swimtime="00:01:14.38" />
                    <SPLIT distance="150" swimtime="00:01:54.68" />
                    <SPLIT distance="200" swimtime="00:02:35.30" />
                    <SPLIT distance="250" swimtime="00:03:16.01" />
                    <SPLIT distance="300" swimtime="00:03:57.30" />
                    <SPLIT distance="350" swimtime="00:04:38.69" />
                    <SPLIT distance="400" swimtime="00:05:20.42" />
                    <SPLIT distance="450" swimtime="00:06:01.77" />
                    <SPLIT distance="500" swimtime="00:06:43.76" />
                    <SPLIT distance="550" swimtime="00:07:24.72" />
                    <SPLIT distance="600" swimtime="00:08:06.45" />
                    <SPLIT distance="650" swimtime="00:08:47.98" />
                    <SPLIT distance="700" swimtime="00:09:28.31" />
                    <SPLIT distance="750" swimtime="00:10:07.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="458" swimtime="00:01:11.68" resultid="11391" heatid="11797" lane="4" entrytime="00:01:11.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 8.5 - Totalmente submerso durante o nado.  (Tempo: 17:56)" eventid="1286" status="DSQ" swimtime="00:03:00.96" resultid="11392" heatid="11813" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                    <SPLIT distance="100" swimtime="00:01:22.13" />
                    <SPLIT distance="150" swimtime="00:02:12.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Pazinato" birthdate="2011-01-05" gender="M" nation="BRA" license="368149" athleteid="11435" externalid="368149">
              <RESULTS>
                <RESULT eventid="1122" points="305" swimtime="00:01:11.73" resultid="11436" heatid="11746" lane="6" entrytime="00:01:13.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="356" swimtime="00:00:28.42" resultid="11437" heatid="11766" lane="6" entrytime="00:00:29.01" entrycourse="SCM" />
                <RESULT eventid="1316" points="358" swimtime="00:01:03.12" resultid="11438" heatid="11835" lane="5" entrytime="00:01:02.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="334" reactiontime="+69" swimtime="00:02:32.15" resultid="11439" heatid="11810" lane="6" entrytime="00:02:48.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                    <SPLIT distance="100" swimtime="00:01:13.24" />
                    <SPLIT distance="150" swimtime="00:01:53.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Dias Rezende" birthdate="2016-03-04" gender="F" nation="BRA" license="406930" athleteid="11533" externalid="406930">
              <RESULTS>
                <RESULT eventid="1178" status="DNS" swimtime="00:00:00.00" resultid="11534" heatid="11768" lane="2" entrytime="00:01:00.32" entrycourse="SCM" />
                <RESULT eventid="1102" status="DNS" swimtime="00:00:00.00" resultid="11535" heatid="11735" lane="5" entrytime="00:01:06.63" entrycourse="SCM" />
                <RESULT eventid="1298" status="DNS" swimtime="00:00:00.00" resultid="11536" heatid="11820" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Guinoza" birthdate="2013-01-06" gender="F" nation="BRA" license="392012" athleteid="11487" externalid="392012">
              <RESULTS>
                <RESULT eventid="1178" points="269" swimtime="00:00:35.48" resultid="11488" heatid="11771" lane="4" entrytime="00:00:37.98" entrycourse="SCM" />
                <RESULT eventid="1102" points="229" swimtime="00:00:46.33" resultid="11489" heatid="11736" lane="3" entrytime="00:00:48.61" entrycourse="SCM" />
                <RESULT eventid="1298" status="DNS" swimtime="00:00:00.00" resultid="11490" heatid="11819" lane="2" />
                <RESULT eventid="1228" points="199" swimtime="00:01:46.71" resultid="11491" heatid="11788" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Correa Mendes" birthdate="2015-05-01" gender="M" nation="BRA" license="422089" athleteid="11554" externalid="422089">
              <RESULTS>
                <RESULT eventid="1183" points="82" swimtime="00:00:46.29" resultid="11555" heatid="11774" lane="1" entrytime="00:00:48.56" entrycourse="SCM" />
                <RESULT eventid="1107" points="94" swimtime="00:00:54.84" resultid="11556" heatid="11737" lane="4" entrytime="00:00:56.87" entrycourse="SCM" />
                <RESULT eventid="1331" points="75" swimtime="00:01:56.54" resultid="11557" heatid="11842" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monique" lastname="Istake" birthdate="2012-04-03" gender="F" nation="BRA" license="372023" athleteid="11406" externalid="372023">
              <RESULTS>
                <RESULT eventid="1142" points="324" swimtime="00:01:18.63" resultid="11407" heatid="11752" lane="5" entrytime="00:01:19.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1162" points="411" swimtime="00:00:30.82" resultid="11408" heatid="11761" lane="6" entrytime="00:00:31.77" entrycourse="SCM" />
                <RESULT comment="SW 8.5 - Totalmente submerso durante o nado.  (Tempo: 17:51)" eventid="1278" status="DSQ" swimtime="00:03:20.45" resultid="11409" heatid="11812" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.02" />
                    <SPLIT distance="150" swimtime="00:02:26.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="355" reactiontime="+153" swimtime="00:05:26.54" resultid="11410" heatid="11780" lane="5" entrytime="00:05:37.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.63" />
                    <SPLIT distance="100" swimtime="00:01:15.51" />
                    <SPLIT distance="150" swimtime="00:01:57.75" />
                    <SPLIT distance="200" swimtime="00:02:40.06" />
                    <SPLIT distance="250" swimtime="00:03:23.00" />
                    <SPLIT distance="300" swimtime="00:04:06.10" />
                    <SPLIT distance="350" swimtime="00:04:47.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Traci Rodrigues" birthdate="2011-03-06" gender="M" nation="BRA" license="406927" athleteid="11398" externalid="406927">
              <RESULTS>
                <RESULT eventid="1170" points="260" swimtime="00:00:31.55" resultid="11399" heatid="11764" lane="1" entrytime="00:00:34.14" entrycourse="SCM" />
                <RESULT eventid="1316" points="259" swimtime="00:01:10.34" resultid="11400" heatid="11833" lane="2" entrytime="00:01:16.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="214" swimtime="00:01:32.28" resultid="11401" heatid="11794" lane="2" entrytime="00:01:39.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Drapzichinski" birthdate="2015-08-21" gender="M" nation="BRA" license="391848" athleteid="11482" externalid="391848">
              <RESULTS>
                <RESULT eventid="1081" points="134" swimtime="00:03:13.80" resultid="11483" heatid="11729" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.18" />
                    <SPLIT distance="100" swimtime="00:01:31.29" />
                    <SPLIT distance="150" swimtime="00:02:25.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="170" swimtime="00:00:36.36" resultid="11484" heatid="11775" lane="4" entrytime="00:00:37.75" entrycourse="SCM" />
                <RESULT eventid="1331" points="124" swimtime="00:01:38.67" resultid="11485" heatid="11843" lane="2" entrytime="00:01:36.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1253" points="122" reactiontime="+83" swimtime="00:00:44.47" resultid="11486" heatid="11802" lane="5" entrytime="00:00:44.82" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Magalhães Rezende" birthdate="2010-05-29" gender="F" nation="BRA" license="366960" athleteid="11416" externalid="366960">
              <RESULTS>
                <RESULT eventid="1060" points="348" swimtime="00:02:36.70" resultid="11417" heatid="11722" lane="3" entrytime="00:02:34.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.75" />
                    <SPLIT distance="100" swimtime="00:01:13.70" />
                    <SPLIT distance="150" swimtime="00:01:54.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="304" swimtime="00:11:49.78" resultid="11418" heatid="11777" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                    <SPLIT distance="100" swimtime="00:01:18.69" />
                    <SPLIT distance="150" swimtime="00:02:02.61" />
                    <SPLIT distance="200" swimtime="00:02:46.70" />
                    <SPLIT distance="250" swimtime="00:03:31.65" />
                    <SPLIT distance="300" swimtime="00:04:16.48" />
                    <SPLIT distance="350" swimtime="00:05:01.89" />
                    <SPLIT distance="400" swimtime="00:05:47.53" />
                    <SPLIT distance="450" swimtime="00:06:33.09" />
                    <SPLIT distance="500" swimtime="00:07:18.72" />
                    <SPLIT distance="550" swimtime="00:08:04.12" />
                    <SPLIT distance="600" swimtime="00:08:50.08" />
                    <SPLIT distance="650" swimtime="00:09:35.45" />
                    <SPLIT distance="700" swimtime="00:10:20.70" />
                    <SPLIT distance="750" swimtime="00:11:05.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1308" points="371" swimtime="00:01:09.92" resultid="11419" heatid="11829" lane="3" entrytime="00:01:10.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="322" swimtime="00:05:37.22" resultid="11420" heatid="11780" lane="2" entrytime="00:05:37.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                    <SPLIT distance="100" swimtime="00:01:16.22" />
                    <SPLIT distance="150" swimtime="00:01:57.81" />
                    <SPLIT distance="200" swimtime="00:02:41.13" />
                    <SPLIT distance="250" swimtime="00:03:25.63" />
                    <SPLIT distance="300" swimtime="00:04:09.79" />
                    <SPLIT distance="350" swimtime="00:04:53.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Catarina" lastname="Benassi Galvani" birthdate="2015-04-20" gender="F" nation="BRA" license="422153" athleteid="11558" externalid="422153">
              <RESULTS>
                <RESULT eventid="1178" points="146" swimtime="00:00:43.54" resultid="11559" heatid="11769" lane="3" entrytime="00:00:49.90" entrycourse="SCM" />
                <RESULT eventid="1102" points="93" swimtime="00:01:02.40" resultid="11560" heatid="11735" lane="6" entrytime="00:01:09.85" entrycourse="SCM" />
                <RESULT eventid="1298" points="118" swimtime="00:01:42.37" resultid="11561" heatid="11820" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18151" nation="BRA" region="PR" clubid="11253" name="Clube Uniao Recreativo Palmense" shortname="Clube União">
          <ATHLETES>
            <ATHLETE firstname="Luiza" lastname="Langaro Spaniol" birthdate="2013-06-18" gender="F" nation="BRA" license="406600" athleteid="11254" externalid="406600">
              <RESULTS>
                <RESULT eventid="1112" points="331" reactiontime="+76" swimtime="00:01:19.29" resultid="11255" heatid="11742" lane="1" entrytime="00:01:15.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="387" swimtime="00:00:31.46" resultid="11256" heatid="11772" lane="2" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1298" points="338" swimtime="00:01:12.09" resultid="11257" heatid="11822" lane="3" entrytime="00:01:08.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="340" swimtime="00:01:29.26" resultid="11258" heatid="11790" lane="3" entrytime="00:01:25.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="36" nation="BRA" region="PR" clubid="11259" name="Associação Atlética Comercial" shortname="Comercial Cascavel">
          <ATHLETES>
            <ATHLETE firstname="Marianna" lastname="Galvao Oliveira" birthdate="2014-03-18" gender="F" nation="BRA" license="390835" athleteid="11324" externalid="390835">
              <RESULTS>
                <RESULT eventid="1112" points="206" reactiontime="+67" swimtime="00:01:32.81" resultid="11325" heatid="11739" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="278" swimtime="00:00:35.11" resultid="11326" heatid="11771" lane="3" entrytime="00:00:37.78" entrycourse="SCM" />
                <RESULT eventid="1228" points="292" swimtime="00:01:33.90" resultid="11327" heatid="11789" lane="4" entrytime="00:01:36.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="260" swimtime="00:03:10.72" resultid="11328" heatid="11844" lane="3" entrytime="00:03:25.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.42" />
                    <SPLIT distance="100" swimtime="00:01:33.89" />
                    <SPLIT distance="150" swimtime="00:02:26.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Larissa" lastname="Yukari Kawai" birthdate="2014-03-13" gender="F" nation="BRA" license="421485" athleteid="11371" externalid="421485">
              <RESULTS>
                <RESULT eventid="1178" points="160" swimtime="00:00:42.22" resultid="11372" heatid="11770" lane="5" entrytime="00:00:44.32" entrycourse="SCM" />
                <RESULT eventid="1102" points="153" swimtime="00:00:53.02" resultid="11373" heatid="11736" lane="1" entrytime="00:00:56.31" entrycourse="SCM" />
                <RESULT eventid="1228" points="180" swimtime="00:01:50.26" resultid="11374" heatid="11788" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.22" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 6.2 - Deixou a posição de costas, exceto ao executar uma virada.  (Tempo: 17:13)" eventid="1248" reactiontime="+101" status="DSQ" swimtime="00:00:46.03" resultid="11375" heatid="11800" lane="5" entrytime="00:00:46.89" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Luis Lottermann" birthdate="2014-10-08" gender="M" nation="BRA" license="382237" athleteid="11289" externalid="382237">
              <RESULTS>
                <RESULT eventid="1152" points="150" swimtime="00:01:29.75" resultid="11290" heatid="11753" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="228" swimtime="00:02:42.61" resultid="11291" heatid="11729" lane="3" entrytime="00:02:42.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                    <SPLIT distance="100" swimtime="00:01:19.13" />
                    <SPLIT distance="150" swimtime="00:02:03.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="191" swimtime="00:03:10.06" resultid="11292" heatid="11846" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.00" />
                    <SPLIT distance="100" swimtime="00:01:29.50" />
                    <SPLIT distance="150" swimtime="00:02:28.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1214" points="199" swimtime="00:06:03.20" resultid="11293" heatid="11782" lane="5" entrytime="00:06:08.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.73" />
                    <SPLIT distance="100" swimtime="00:01:27.46" />
                    <SPLIT distance="150" swimtime="00:02:13.69" />
                    <SPLIT distance="200" swimtime="00:03:00.67" />
                    <SPLIT distance="250" swimtime="00:03:49.26" />
                    <SPLIT distance="300" swimtime="00:04:36.47" />
                    <SPLIT distance="350" swimtime="00:05:23.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Flavia" lastname="De Metz" birthdate="2011-01-07" gender="F" nation="BRA" license="390846" athleteid="11334" externalid="390846">
              <RESULTS>
                <RESULT eventid="1112" points="337" reactiontime="+73" swimtime="00:01:18.87" resultid="11335" heatid="11742" lane="6" entrytime="00:01:18.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1262" points="370" reactiontime="+79" swimtime="00:02:45.66" resultid="11336" heatid="11808" lane="2" entrytime="00:02:44.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.94" />
                    <SPLIT distance="100" swimtime="00:01:21.13" />
                    <SPLIT distance="150" swimtime="00:02:04.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="370" swimtime="00:02:49.69" resultid="11337" heatid="11845" lane="2" entrytime="00:02:53.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                    <SPLIT distance="100" swimtime="00:01:19.65" />
                    <SPLIT distance="150" swimtime="00:02:12.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Claudio" lastname="Rohnelt" birthdate="2010-03-08" gender="M" nation="BRA" license="357954" athleteid="11260" externalid="357954">
              <RESULTS>
                <RESULT eventid="1152" points="343" swimtime="00:01:08.24" resultid="11261" heatid="11757" lane="1" entrytime="00:01:09.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="362" swimtime="00:02:19.40" resultid="11262" heatid="11725" lane="5" entrytime="00:02:17.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                    <SPLIT distance="100" swimtime="00:01:07.02" />
                    <SPLIT distance="150" swimtime="00:01:43.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="331" swimtime="00:02:34.41" resultid="11263" heatid="11815" lane="6" entrytime="00:02:36.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                    <SPLIT distance="100" swimtime="00:01:14.62" />
                    <SPLIT distance="150" swimtime="00:01:54.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="371" swimtime="00:02:32.50" resultid="11264" heatid="11849" lane="3" entrytime="00:02:35.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                    <SPLIT distance="100" swimtime="00:01:12.44" />
                    <SPLIT distance="150" swimtime="00:01:57.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raul" lastname="Bonamigo" birthdate="2010-12-01" gender="M" nation="BRA" license="344397" athleteid="11304" externalid="344397">
              <RESULTS>
                <RESULT eventid="1152" points="318" swimtime="00:01:09.96" resultid="11305" heatid="11757" lane="5" entrytime="00:01:08.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="473" swimtime="00:02:07.45" resultid="11306" heatid="11725" lane="3" entrytime="00:02:11.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.84" />
                    <SPLIT distance="100" swimtime="00:01:00.37" />
                    <SPLIT distance="150" swimtime="00:01:33.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="438" swimtime="00:02:24.31" resultid="11307" heatid="11850" lane="5" entrytime="00:02:25.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.26" />
                    <SPLIT distance="100" swimtime="00:01:07.80" />
                    <SPLIT distance="150" swimtime="00:01:51.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1214" points="477" swimtime="00:04:31.52" resultid="11308" heatid="11783" lane="4" entrytime="00:04:31.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                    <SPLIT distance="100" swimtime="00:01:04.27" />
                    <SPLIT distance="150" swimtime="00:01:38.28" />
                    <SPLIT distance="200" swimtime="00:02:12.57" />
                    <SPLIT distance="250" swimtime="00:02:47.18" />
                    <SPLIT distance="300" swimtime="00:03:21.84" />
                    <SPLIT distance="350" swimtime="00:03:57.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Breno" lastname="Zanella Janke" birthdate="2011-04-26" gender="M" nation="BRA" license="365697" athleteid="11270" externalid="365697">
              <RESULTS>
                <RESULT eventid="1152" points="342" swimtime="00:01:08.26" resultid="11271" heatid="11757" lane="4" entrytime="00:01:07.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1094" points="354" swimtime="00:02:49.83" resultid="11272" heatid="11733" lane="6" entrytime="00:02:50.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.62" />
                    <SPLIT distance="100" swimtime="00:01:20.39" />
                    <SPLIT distance="150" swimtime="00:02:05.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="387" swimtime="00:01:15.84" resultid="11273" heatid="11796" lane="4" entrytime="00:01:18.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="327" swimtime="00:02:35.09" resultid="11274" heatid="11814" lane="3" entrytime="00:02:42.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                    <SPLIT distance="100" swimtime="00:01:13.20" />
                    <SPLIT distance="150" swimtime="00:01:54.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="Gabriel Dalchau" birthdate="2014-08-27" gender="M" nation="BRA" license="402118" athleteid="11348" externalid="402118">
              <RESULTS>
                <RESULT eventid="1122" points="141" swimtime="00:01:32.66" resultid="11349" heatid="11744" lane="2" entrytime="00:01:31.46" entrycourse="SCM" />
                <RESULT eventid="1081" points="157" swimtime="00:03:03.89" resultid="11350" heatid="11728" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.03" />
                    <SPLIT distance="100" swimtime="00:01:27.36" />
                    <SPLIT distance="150" swimtime="00:02:16.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="145" swimtime="00:03:28.63" resultid="11351" heatid="11847" lane="3" entrytime="00:03:23.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.84" />
                    <SPLIT distance="100" swimtime="00:01:42.26" />
                    <SPLIT distance="150" swimtime="00:02:43.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1214" points="153" swimtime="00:06:36.30" resultid="11352" heatid="11782" lane="6" entrytime="00:06:28.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.69" />
                    <SPLIT distance="100" swimtime="00:01:33.29" />
                    <SPLIT distance="150" swimtime="00:02:23.79" />
                    <SPLIT distance="200" swimtime="00:03:15.99" />
                    <SPLIT distance="250" swimtime="00:04:07.89" />
                    <SPLIT distance="300" swimtime="00:04:58.93" />
                    <SPLIT distance="350" swimtime="00:05:50.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Cordeiro Silva" birthdate="2011-09-04" gender="M" nation="BRA" license="380664" athleteid="11284" externalid="380664">
              <RESULTS>
                <RESULT eventid="1152" points="214" swimtime="00:01:19.77" resultid="11285" heatid="11754" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1094" points="356" swimtime="00:02:49.45" resultid="11286" heatid="11732" lane="3" entrytime="00:02:55.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.88" />
                    <SPLIT distance="100" swimtime="00:01:22.08" />
                    <SPLIT distance="150" swimtime="00:02:04.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="342" swimtime="00:01:19.04" resultid="11287" heatid="11796" lane="5" entrytime="00:01:23.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="306" swimtime="00:02:42.67" resultid="11288" heatid="11849" lane="1" entrytime="00:02:48.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                    <SPLIT distance="100" swimtime="00:01:22.84" />
                    <SPLIT distance="150" swimtime="00:02:04.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Bonamigo" birthdate="2013-06-25" gender="M" nation="BRA" license="365484" athleteid="11319" externalid="365484">
              <RESULTS>
                <RESULT eventid="1107" points="222" swimtime="00:00:41.19" resultid="11320" heatid="11738" lane="3" entrytime="00:00:39.46" entrycourse="SCM" />
                <RESULT eventid="1137" points="220" swimtime="00:00:36.00" resultid="11321" heatid="11749" lane="3" entrytime="00:00:36.18" entrycourse="SCM" />
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente., Na volta dos 75m." eventid="1238" status="DSQ" swimtime="00:01:29.10" resultid="11322" heatid="11795" lane="4" entrytime="00:01:28.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="251" swimtime="00:02:53.57" resultid="11323" heatid="11849" lane="6" entrytime="00:02:51.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                    <SPLIT distance="100" swimtime="00:01:25.37" />
                    <SPLIT distance="150" swimtime="00:02:14.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanna" lastname="Bertelli Weirich" birthdate="2011-03-18" gender="F" nation="BRA" license="369534" athleteid="11275" externalid="369534">
              <RESULTS>
                <RESULT eventid="1142" points="338" swimtime="00:01:17.53" resultid="11276" heatid="11752" lane="4" entrytime="00:01:13.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="395" swimtime="00:02:30.22" resultid="11277" heatid="11723" lane="5" entrytime="00:02:22.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.15" />
                    <SPLIT distance="100" swimtime="00:01:11.32" />
                    <SPLIT distance="150" swimtime="00:01:50.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="382" swimtime="00:02:44.71" resultid="11278" heatid="11812" lane="3" entrytime="00:02:41.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.60" />
                    <SPLIT distance="100" swimtime="00:01:18.27" />
                    <SPLIT distance="150" swimtime="00:02:00.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benicio" lastname="Hermisdorff Bruning" birthdate="2015-06-22" gender="M" nation="BRA" license="414000" athleteid="11363" externalid="414000">
              <RESULTS>
                <RESULT eventid="1331" points="122" swimtime="00:01:39.34" resultid="11364" heatid="11843" lane="5" entrytime="00:01:42.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1253" points="130" reactiontime="+60" swimtime="00:00:43.55" resultid="11365" heatid="11802" lane="1" entrytime="00:00:46.57" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Pedro Serafini" birthdate="2012-05-15" gender="M" nation="BRA" license="365488" athleteid="11314" externalid="365488">
              <RESULTS>
                <RESULT eventid="1152" points="239" swimtime="00:01:16.91" resultid="11315" heatid="11756" lane="1" entrytime="00:01:24.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="359" swimtime="00:10:19.23" resultid="11316" heatid="11778" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.46" />
                    <SPLIT distance="100" swimtime="00:01:14.10" />
                    <SPLIT distance="150" swimtime="00:01:52.90" />
                    <SPLIT distance="200" swimtime="00:02:32.32" />
                    <SPLIT distance="250" swimtime="00:03:11.74" />
                    <SPLIT distance="300" swimtime="00:03:50.75" />
                    <SPLIT distance="350" swimtime="00:04:30.46" />
                    <SPLIT distance="400" swimtime="00:05:10.24" />
                    <SPLIT distance="450" swimtime="00:05:49.57" />
                    <SPLIT distance="500" swimtime="00:06:29.26" />
                    <SPLIT distance="550" swimtime="00:07:08.43" />
                    <SPLIT distance="600" swimtime="00:07:47.07" />
                    <SPLIT distance="650" swimtime="00:08:25.90" />
                    <SPLIT distance="700" swimtime="00:09:04.52" />
                    <SPLIT distance="750" swimtime="00:09:43.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="285" swimtime="00:02:46.44" resultid="11317" heatid="11848" lane="3" entrytime="00:02:52.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.71" />
                    <SPLIT distance="100" swimtime="00:01:21.73" />
                    <SPLIT distance="150" swimtime="00:02:09.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1214" points="364" swimtime="00:04:57.05" resultid="11318" heatid="11782" lane="3" entrytime="00:05:07.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                    <SPLIT distance="100" swimtime="00:01:11.06" />
                    <SPLIT distance="150" swimtime="00:01:49.00" />
                    <SPLIT distance="200" swimtime="00:02:27.29" />
                    <SPLIT distance="250" swimtime="00:03:05.58" />
                    <SPLIT distance="300" swimtime="00:03:43.88" />
                    <SPLIT distance="350" swimtime="00:04:21.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="Menegazzi Daga" birthdate="2014-12-05" gender="M" nation="BRA" license="414003" athleteid="11366" externalid="414003">
              <RESULTS>
                <RESULT eventid="1122" points="92" reactiontime="+86" swimtime="00:01:46.78" resultid="11367" heatid="11743" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="66" swimtime="00:00:49.88" resultid="11368" heatid="11774" lane="4" entrytime="00:00:45.23" entrycourse="SCM" />
                <RESULT eventid="1238" points="113" swimtime="00:01:54.32" resultid="11369" heatid="11793" lane="2" entrytime="00:02:06.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="114" swimtime="00:03:45.64" resultid="11370" heatid="11847" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.51" />
                    <SPLIT distance="100" swimtime="00:01:49.08" />
                    <SPLIT distance="150" swimtime="00:02:51.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexia" lastname="Moura Ticianelli" birthdate="2013-04-04" gender="F" nation="BRA" license="406785" athleteid="11376" externalid="406785">
              <RESULTS>
                <RESULT eventid="1112" points="305" reactiontime="+70" swimtime="00:01:21.51" resultid="11377" heatid="11741" lane="5" entrytime="00:01:22.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="322" swimtime="00:00:33.42" resultid="11378" heatid="11772" lane="1" entrytime="00:00:34.95" entrycourse="SCM" />
                <RESULT eventid="1334" points="317" swimtime="00:02:58.62" resultid="11379" heatid="11845" lane="1" entrytime="00:03:01.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.59" />
                    <SPLIT distance="100" swimtime="00:01:24.05" />
                    <SPLIT distance="150" swimtime="00:02:18.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="306" reactiontime="+72" swimtime="00:00:37.43" resultid="11380" heatid="11800" lane="3" entrytime="00:00:38.99" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Assakura" birthdate="2010-06-29" gender="F" nation="BRA" license="376473" athleteid="11299" externalid="376473">
              <RESULTS>
                <RESULT eventid="1142" points="334" swimtime="00:01:17.89" resultid="11300" heatid="11751" lane="4" entrytime="00:01:24.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1086" points="494" swimtime="00:02:50.20" resultid="11301" heatid="11731" lane="3" entrytime="00:02:48.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                    <SPLIT distance="100" swimtime="00:01:22.20" />
                    <SPLIT distance="150" swimtime="00:02:07.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="439" swimtime="00:01:22.02" resultid="11302" heatid="11791" lane="1" entrytime="00:01:20.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="486" swimtime="00:04:54.17" resultid="11303" heatid="11779" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                    <SPLIT distance="100" swimtime="00:01:08.81" />
                    <SPLIT distance="150" swimtime="00:01:45.89" />
                    <SPLIT distance="200" swimtime="00:02:23.40" />
                    <SPLIT distance="250" swimtime="00:03:01.75" />
                    <SPLIT distance="300" swimtime="00:03:39.89" />
                    <SPLIT distance="350" swimtime="00:04:17.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="Bortoli Da Silva" birthdate="2010-09-30" gender="M" nation="BRA" license="365500" athleteid="11358" externalid="365500">
              <RESULTS>
                <RESULT eventid="1152" points="327" swimtime="00:01:09.32" resultid="11359" heatid="11756" lane="3" entrytime="00:01:10.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="379" swimtime="00:02:17.23" resultid="11360" heatid="11725" lane="4" entrytime="00:02:15.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.27" />
                    <SPLIT distance="100" swimtime="00:01:06.26" />
                    <SPLIT distance="150" swimtime="00:01:42.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="327" swimtime="00:02:34.99" resultid="11361" heatid="11814" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                    <SPLIT distance="100" swimtime="00:01:12.01" />
                    <SPLIT distance="150" swimtime="00:01:52.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="365" swimtime="00:02:33.30" resultid="11362" heatid="11849" lane="4" entrytime="00:02:35.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:16.22" />
                    <SPLIT distance="150" swimtime="00:01:59.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Macedo Medeiros" birthdate="2012-05-12" gender="M" nation="BRA" license="392015" athleteid="11343" externalid="392015">
              <RESULTS>
                <RESULT eventid="1152" points="151" swimtime="00:01:29.61" resultid="11344" heatid="11755" lane="5" entrytime="00:01:37.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1094" points="244" swimtime="00:03:12.07" resultid="11345" heatid="11732" lane="2" entrytime="00:03:20.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.87" />
                    <SPLIT distance="100" swimtime="00:01:32.90" />
                    <SPLIT distance="150" swimtime="00:02:23.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="228" swimtime="00:01:30.44" resultid="11346" heatid="11795" lane="1" entrytime="00:01:34.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="226" swimtime="00:02:59.98" resultid="11347" heatid="11848" lane="1" entrytime="00:03:03.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.95" />
                    <SPLIT distance="100" swimtime="00:01:32.25" />
                    <SPLIT distance="150" swimtime="00:02:21.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Ramirez Vasconcelos" birthdate="2011-04-06" gender="M" nation="BRA" license="392013" athleteid="11338" externalid="392013">
              <RESULTS>
                <RESULT eventid="1152" points="325" swimtime="00:01:09.48" resultid="11339" heatid="11756" lane="4" entrytime="00:01:11.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="400" swimtime="00:02:14.78" resultid="11340" heatid="11725" lane="2" entrytime="00:02:16.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                    <SPLIT distance="100" swimtime="00:01:03.88" />
                    <SPLIT distance="150" swimtime="00:01:39.01" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 6.2 - Deixou a posição de costas, exceto ao executar uma virada.  (Tempo: 19:59), Na volta dos 100m (Costas, Medley Individual)." eventid="1344" status="DSQ" swimtime="00:02:32.08" resultid="11341" heatid="11850" lane="6" entrytime="00:02:32.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                    <SPLIT distance="100" swimtime="00:01:13.02" />
                    <SPLIT distance="150" swimtime="00:01:56.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1214" points="412" swimtime="00:04:45.05" resultid="11342" heatid="11782" lane="4" entrytime="00:05:10.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.79" />
                    <SPLIT distance="100" swimtime="00:01:05.95" />
                    <SPLIT distance="150" swimtime="00:01:42.72" />
                    <SPLIT distance="200" swimtime="00:02:19.53" />
                    <SPLIT distance="250" swimtime="00:02:56.53" />
                    <SPLIT distance="300" swimtime="00:03:33.77" />
                    <SPLIT distance="350" swimtime="00:04:09.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="11888" points="407" swimtime="00:05:16.60" resultid="11899" heatid="11898" lane="1" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                    <SPLIT distance="100" swimtime="00:01:12.06" />
                    <SPLIT distance="150" swimtime="00:01:53.55" />
                    <SPLIT distance="200" swimtime="00:02:36.82" />
                    <SPLIT distance="250" swimtime="00:03:17.88" />
                    <SPLIT distance="300" swimtime="00:04:02.56" />
                    <SPLIT distance="350" swimtime="00:04:40.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Luisa Lottermann" birthdate="2011-08-26" gender="F" nation="BRA" license="382238" athleteid="11294" externalid="382238">
              <RESULTS>
                <RESULT eventid="1142" points="214" swimtime="00:01:30.23" resultid="11295" heatid="11751" lane="5" entrytime="00:01:27.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1086" points="402" swimtime="00:03:02.27" resultid="11296" heatid="11731" lane="2" entrytime="00:02:59.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.65" />
                    <SPLIT distance="100" swimtime="00:01:28.09" />
                    <SPLIT distance="150" swimtime="00:02:15.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="373" swimtime="00:01:26.63" resultid="11297" heatid="11791" lane="6" entrytime="00:01:25.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="248" swimtime="00:03:10.14" resultid="11298" heatid="11812" lane="2" entrytime="00:03:07.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.96" />
                    <SPLIT distance="100" swimtime="00:01:32.86" />
                    <SPLIT distance="150" swimtime="00:02:21.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Emanuel Rech" birthdate="2013-12-02" gender="M" nation="BRA" license="380660" athleteid="11279" externalid="380660">
              <RESULTS>
                <RESULT eventid="1122" points="220" swimtime="00:01:19.98" resultid="11280" heatid="11745" lane="1" entrytime="00:01:23.04" entrycourse="SCM" />
                <RESULT eventid="1183" points="266" swimtime="00:00:31.32" resultid="11281" heatid="11776" lane="2" entrytime="00:00:33.26" entrycourse="SCM" />
                <RESULT eventid="1344" points="242" swimtime="00:02:55.90" resultid="11282" heatid="11848" lane="5" entrytime="00:03:00.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.64" />
                    <SPLIT distance="150" swimtime="00:02:18.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1253" points="215" reactiontime="+61" swimtime="00:00:36.89" resultid="11283" heatid="11802" lane="3" entrytime="00:00:37.23" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laisa" lastname="Bernardini" birthdate="2012-06-25" gender="F" nation="BRA" license="390843" athleteid="11329" externalid="390843">
              <RESULTS>
                <RESULT eventid="1142" points="204" swimtime="00:01:31.67" resultid="11330" heatid="11751" lane="6" entrytime="00:01:37.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1086" points="314" swimtime="00:03:17.95" resultid="11331" heatid="11730" lane="4" entrytime="00:03:27.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.24" />
                    <SPLIT distance="100" swimtime="00:01:37.44" />
                    <SPLIT distance="150" swimtime="00:02:28.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="297" swimtime="00:01:33.45" resultid="11332" heatid="11789" lane="3" entrytime="00:01:36.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="321" swimtime="00:02:57.82" resultid="11333" heatid="11845" lane="5" entrytime="00:03:01.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.76" />
                    <SPLIT distance="100" swimtime="00:01:28.57" />
                    <SPLIT distance="150" swimtime="00:02:18.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Alves Serafini" birthdate="2008-04-15" gender="M" nation="BRA" license="351644" athleteid="11309" externalid="351644">
              <RESULTS>
                <RESULT eventid="1152" points="445" swimtime="00:01:02.55" resultid="11310" heatid="11758" lane="2" entrytime="00:01:00.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="445" swimtime="00:02:10.07" resultid="11311" heatid="11726" lane="5" entrytime="00:02:04.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                    <SPLIT distance="100" swimtime="00:01:00.81" />
                    <SPLIT distance="150" swimtime="00:01:35.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="477" swimtime="00:02:16.68" resultid="11312" heatid="11815" lane="3" entrytime="00:02:14.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                    <SPLIT distance="100" swimtime="00:01:04.98" />
                    <SPLIT distance="150" swimtime="00:01:38.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1214" points="520" swimtime="00:04:23.89" resultid="11313" heatid="11783" lane="3" entrytime="00:04:24.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.18" />
                    <SPLIT distance="100" swimtime="00:01:02.59" />
                    <SPLIT distance="150" swimtime="00:01:35.43" />
                    <SPLIT distance="200" swimtime="00:02:08.49" />
                    <SPLIT distance="250" swimtime="00:02:41.94" />
                    <SPLIT distance="300" swimtime="00:03:15.87" />
                    <SPLIT distance="350" swimtime="00:03:50.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Vieira Rohnelt" birthdate="2012-05-03" gender="M" nation="BRA" license="365692" athleteid="11265" externalid="365692">
              <RESULTS>
                <RESULT eventid="1122" points="202" swimtime="00:01:22.33" resultid="11266" heatid="11745" lane="5" entrytime="00:01:22.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="269" swimtime="00:02:33.88" resultid="11267" heatid="11724" lane="4" entrytime="00:02:45.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                    <SPLIT distance="100" swimtime="00:01:13.54" />
                    <SPLIT distance="150" swimtime="00:01:54.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="230" reactiontime="+85" swimtime="00:02:52.23" resultid="11268" heatid="11809" lane="2" entrytime="00:02:56.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.05" />
                    <SPLIT distance="100" swimtime="00:01:24.86" />
                    <SPLIT distance="150" swimtime="00:02:08.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="243" swimtime="00:02:55.60" resultid="11269" heatid="11848" lane="4" entrytime="00:02:56.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.22" />
                    <SPLIT distance="100" swimtime="00:01:26.56" />
                    <SPLIT distance="150" swimtime="00:02:17.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Henrique Marca Dos Santos" birthdate="2015-03-28" gender="M" nation="BRA" license="406695" athleteid="11353" externalid="406695">
              <RESULTS>
                <RESULT eventid="1183" points="190" swimtime="00:00:35.05" resultid="11354" heatid="11776" lane="6" entrytime="00:00:36.12" entrycourse="SCM" />
                <RESULT eventid="1107" points="149" swimtime="00:00:46.97" resultid="11355" heatid="11738" lane="5" entrytime="00:00:53.14" entrycourse="SCM" />
                <RESULT eventid="1331" points="191" swimtime="00:01:25.46" resultid="11356" heatid="11843" lane="3" entrytime="00:01:31.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="225" swimtime="00:01:13.69" resultid="11357" heatid="11826" lane="4" entrytime="00:01:16.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="1035" nation="BRA" region="PR" clubid="11574" name="Fundação De Esportes De Campo Mourão" shortname="Fecam">
          <ATHLETES>
            <ATHLETE firstname="Fabricio" lastname="Campos Faria" birthdate="2013-09-15" gender="M" nation="BRA" license="422156" athleteid="11667" externalid="422156">
              <RESULTS>
                <RESULT eventid="1183" points="177" swimtime="00:00:35.89" resultid="11668" heatid="11775" lane="5" entrytime="00:00:38.28" entrycourse="SCM" />
                <RESULT eventid="1303" status="DNS" swimtime="00:00:00.00" resultid="11669" heatid="11823" lane="3" />
                <RESULT eventid="1253" points="91" reactiontime="+71" swimtime="00:00:49.12" resultid="11670" heatid="11801" lane="4" entrytime="00:00:54.04" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Franca Rebollo" birthdate="2012-09-26" gender="M" nation="BRA" license="385780" athleteid="11575" externalid="385780">
              <RESULTS>
                <RESULT eventid="1122" points="134" swimtime="00:01:34.42" resultid="11576" heatid="11744" lane="1" entrytime="00:01:36.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="155" swimtime="00:00:37.46" resultid="11577" heatid="11763" lane="5" entrytime="00:00:38.24" entrycourse="SCM" />
                <RESULT eventid="1316" points="141" swimtime="00:01:26.06" resultid="11578" heatid="11832" lane="4" entrytime="00:01:25.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="133" reactiontime="+85" swimtime="00:03:26.68" resultid="11579" heatid="11809" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.96" />
                    <SPLIT distance="100" swimtime="00:01:43.61" />
                    <SPLIT distance="150" swimtime="00:02:37.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduarda" lastname="Daleffe Pepino" birthdate="2000-07-09" gender="F" nation="BRA" license="185817" athleteid="11588" externalid="185817">
              <RESULTS>
                <RESULT eventid="1112" points="277" reactiontime="+59" swimtime="00:01:24.17" resultid="11589" heatid="11741" lane="4" entrytime="00:01:22.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1162" points="388" swimtime="00:00:31.42" resultid="11590" heatid="11761" lane="1" entrytime="00:00:31.65" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonia" lastname="Giglini Zambon" birthdate="2015-05-25" gender="F" nation="BRA" license="422157" athleteid="11671" externalid="422157">
              <RESULTS>
                <RESULT eventid="1178" points="102" swimtime="00:00:48.99" resultid="11672" heatid="11769" lane="2" entrytime="00:00:51.66" entrycourse="SCM" />
                <RESULT eventid="1298" points="82" swimtime="00:01:55.34" resultid="11673" heatid="11819" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="67" reactiontime="+61" swimtime="00:01:02.08" resultid="11674" heatid="11798" lane="2" entrytime="00:01:13.44" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Ferreira Batista" birthdate="2012-03-29" gender="F" nation="BRA" license="385779" athleteid="11617" externalid="385779">
              <RESULTS>
                <RESULT eventid="1112" points="223" reactiontime="+65" swimtime="00:01:30.48" resultid="11618" heatid="11740" lane="2" entrytime="00:01:28.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="233" swimtime="00:02:59.14" resultid="11619" heatid="11722" lane="4" entrytime="00:03:00.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                    <SPLIT distance="100" swimtime="00:01:26.08" />
                    <SPLIT distance="150" swimtime="00:02:14.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1162" points="281" swimtime="00:00:34.99" resultid="11620" heatid="11760" lane="1" entrytime="00:00:34.46" entrycourse="SCM" />
                <RESULT eventid="1308" status="DNS" swimtime="00:00:00.00" resultid="11621" heatid="11828" lane="4" entrytime="00:01:18.45" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur" lastname="Setsuo Iechika" birthdate="2013-03-10" gender="M" nation="BRA" license="422155" athleteid="11663" externalid="422155">
              <RESULTS>
                <RESULT eventid="1183" points="103" swimtime="00:00:42.91" resultid="11664" heatid="11774" lane="2" entrytime="00:00:45.74" entrycourse="SCM" />
                <RESULT eventid="1303" points="88" swimtime="00:01:40.59" resultid="11665" heatid="11824" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1253" points="76" reactiontime="+69" swimtime="00:00:52.07" resultid="11666" heatid="11801" lane="3" entrytime="00:00:52.39" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henry" lastname="Sadao Da Silva" birthdate="2012-10-02" gender="M" nation="BRA" license="413907" athleteid="11647" externalid="413907">
              <RESULTS>
                <RESULT eventid="1122" points="108" swimtime="00:01:41.26" resultid="11648" heatid="11744" lane="6" entrytime="00:01:51.97" entrycourse="SCM" />
                <RESULT eventid="1170" points="161" swimtime="00:00:37.00" resultid="11649" heatid="11762" lane="3" entrytime="00:00:43.10" entrycourse="SCM" />
                <RESULT eventid="1316" points="143" swimtime="00:01:25.71" resultid="11650" heatid="11832" lane="6" entrytime="00:01:31.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="112" swimtime="00:03:47.14" resultid="11651" heatid="11846" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.93" />
                    <SPLIT distance="100" swimtime="00:01:48.89" />
                    <SPLIT distance="150" swimtime="00:02:56.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Franco Santos" birthdate="2002-01-03" gender="M" nation="BRA" license="290441" athleteid="11599" externalid="290441">
              <RESULTS>
                <RESULT eventid="1152" points="412" swimtime="00:01:04.16" resultid="11600" heatid="11754" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="535" swimtime="00:00:24.82" resultid="11601" heatid="11767" lane="4" entrytime="00:00:24.83" entrycourse="SCM" />
                <RESULT eventid="1316" points="452" swimtime="00:00:58.39" resultid="11602" heatid="11836" lane="1" entrytime="00:00:56.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.41" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 6.5 - Não terminou a prova enquanto estava de costas.&#10;&#10;&#10;&#10;&#10;&#10;&#10;  (Tempo: 19:59), Na volta dos 100m (Costas, Medley Individual)." eventid="1344" status="DSQ" swimtime="00:02:43.24" resultid="11603" heatid="11850" lane="1" entrytime="00:02:30.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                    <SPLIT distance="100" swimtime="00:01:12.09" />
                    <SPLIT distance="150" swimtime="00:02:04.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaue" lastname="Guilherme Chagas" birthdate="2005-06-29" gender="M" nation="BRA" license="378464" athleteid="11613" externalid="378464">
              <RESULTS>
                <RESULT eventid="1170" points="334" swimtime="00:00:29.05" resultid="11614" heatid="11766" lane="5" entrytime="00:00:28.54" entrycourse="SCM" />
                <RESULT eventid="1316" points="313" swimtime="00:01:06.03" resultid="11615" heatid="11835" lane="2" entrytime="00:01:02.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="251" swimtime="00:01:27.60" resultid="11616" heatid="11796" lane="6" entrytime="00:01:26.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Paulo Pedroso" birthdate="1995-11-14" gender="M" nation="BRA" license="115711" athleteid="11580" externalid="115711">
              <RESULTS>
                <RESULT eventid="1122" points="333" swimtime="00:01:09.71" resultid="11581" heatid="11746" lane="2" entrytime="00:01:09.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="409" swimtime="00:00:27.14" resultid="11582" heatid="11767" lane="1" entrytime="00:00:27.25" entrycourse="SCM" />
                <RESULT eventid="1270" points="288" reactiontime="+61" swimtime="00:02:39.95" resultid="11583" heatid="11810" lane="1" entrytime="00:02:38.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                    <SPLIT distance="150" swimtime="00:01:58.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Keirrison" lastname="Leite Silva" birthdate="2011-08-02" gender="M" nation="BRA" license="392161" athleteid="11591" externalid="392161">
              <RESULTS>
                <RESULT eventid="1170" points="173" swimtime="00:00:36.14" resultid="11592" heatid="11763" lane="4" entrytime="00:00:37.90" entrycourse="SCM" />
                <RESULT eventid="1316" points="157" swimtime="00:01:22.95" resultid="11593" heatid="11832" lane="5" entrytime="00:01:29.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.43" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.4 - Movimentos das pernas não simultâneos.  (Tempo: 16:51), Após a volta dos 50m." eventid="1238" status="DSQ" swimtime="00:01:44.71" resultid="11594" heatid="11793" lane="3" entrytime="00:01:57.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raul" lastname="Massuda Santos" birthdate="2017-10-28" gender="M" nation="BRA" license="424520" athleteid="11685" externalid="424520">
              <RESULTS>
                <RESULT eventid="1326" points="71" swimtime="00:00:48.49" resultid="11686" heatid="11839" lane="4" />
                <RESULT eventid="1260" points="66" swimtime="00:00:25.36" resultid="11687" heatid="11805" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Stipp Silva" birthdate="2009-12-02" gender="M" nation="BRA" license="378462" athleteid="11608" externalid="378462">
              <RESULTS>
                <RESULT eventid="1170" points="463" swimtime="00:00:26.05" resultid="11609" heatid="11767" lane="2" entrytime="00:00:25.94" entrycourse="SCM" />
                <RESULT eventid="1316" points="463" swimtime="00:00:57.96" resultid="11610" heatid="11836" lane="6" entrytime="00:00:57.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="393" swimtime="00:01:15.44" resultid="11611" heatid="11797" lane="1" entrytime="00:01:14.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="374" swimtime="00:02:32.08" resultid="11612" heatid="11846" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                    <SPLIT distance="100" swimtime="00:01:11.58" />
                    <SPLIT distance="150" swimtime="00:01:55.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Capel Adelino" birthdate="2009-04-24" gender="M" nation="BRA" license="422154" athleteid="11660" externalid="422154">
              <RESULTS>
                <RESULT eventid="1170" points="225" swimtime="00:00:33.14" resultid="11661" heatid="11764" lane="2" entrytime="00:00:33.06" entrycourse="SCM" />
                <RESULT eventid="1316" points="191" swimtime="00:01:17.78" resultid="11662" heatid="11832" lane="3" entrytime="00:01:21.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Eduardo Schork Filho" birthdate="2012-12-28" gender="M" nation="BRA" license="413906" athleteid="11643" externalid="413906">
              <RESULTS>
                <RESULT eventid="1170" points="157" swimtime="00:00:37.33" resultid="11644" heatid="11763" lane="2" entrytime="00:00:38.01" entrycourse="SCM" />
                <RESULT eventid="1316" points="125" swimtime="00:01:29.48" resultid="11645" heatid="11832" lane="2" entrytime="00:01:28.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="144" swimtime="00:01:45.25" resultid="11646" heatid="11794" lane="1" entrytime="00:01:49.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Batinga Ponchielli" birthdate="2007-01-18" gender="M" nation="BRA" license="378461" athleteid="11604" externalid="378461">
              <RESULTS>
                <RESULT eventid="1122" points="253" swimtime="00:01:16.36" resultid="11605" heatid="11745" lane="3" entrytime="00:01:14.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="325" swimtime="00:00:29.31" resultid="11606" heatid="11766" lane="1" entrytime="00:00:28.90" entrycourse="SCM" />
                <RESULT eventid="1270" points="208" reactiontime="+76" swimtime="00:02:58.09" resultid="11607" heatid="11809" lane="3" entrytime="00:02:52.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.99" />
                    <SPLIT distance="100" swimtime="00:01:25.09" />
                    <SPLIT distance="150" swimtime="00:02:13.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juliana" lastname="De Oliveira Palo Machado" birthdate="1983-09-28" gender="F" nation="BRA" license="419883" athleteid="11682" externalid="419883">
              <RESULTS>
                <RESULT eventid="1162" points="318" swimtime="00:00:33.56" resultid="11683" heatid="11759" lane="1" />
                <RESULT eventid="1308" status="DNS" swimtime="00:00:00.00" resultid="11684" heatid="11827" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Felipe Damha" birthdate="1987-01-02" gender="M" nation="BRA" license="053982" athleteid="11679" externalid="053982">
              <RESULTS>
                <RESULT eventid="1170" points="456" swimtime="00:00:26.19" resultid="11680" heatid="11762" lane="5" />
                <RESULT eventid="1270" points="314" reactiontime="+81" swimtime="00:02:35.32" resultid="11681" heatid="11810" lane="2" entrytime="00:02:34.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                    <SPLIT distance="100" swimtime="00:01:15.41" />
                    <SPLIT distance="150" swimtime="00:01:54.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Pedroso Silverio" birthdate="1994-11-21" gender="M" nation="BRA" license="115715" athleteid="11584" externalid="115715">
              <RESULTS>
                <RESULT eventid="1196" points="314" swimtime="00:10:47.58" resultid="11585" heatid="11778" lane="4" entrytime="00:10:30.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:13.22" />
                    <SPLIT distance="150" swimtime="00:01:52.20" />
                    <SPLIT distance="200" swimtime="00:02:31.33" />
                    <SPLIT distance="250" swimtime="00:03:11.18" />
                    <SPLIT distance="300" swimtime="00:03:51.24" />
                    <SPLIT distance="350" swimtime="00:04:31.67" />
                    <SPLIT distance="400" swimtime="00:05:12.72" />
                    <SPLIT distance="450" swimtime="00:05:54.28" />
                    <SPLIT distance="500" swimtime="00:06:35.78" />
                    <SPLIT distance="550" swimtime="00:07:17.94" />
                    <SPLIT distance="600" swimtime="00:08:00.12" />
                    <SPLIT distance="650" swimtime="00:08:41.95" />
                    <SPLIT distance="700" swimtime="00:09:24.29" />
                    <SPLIT distance="750" swimtime="00:10:06.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="263" swimtime="00:02:46.74" resultid="11586" heatid="11813" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.08" />
                    <SPLIT distance="100" swimtime="00:01:22.61" />
                    <SPLIT distance="150" swimtime="00:02:06.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1214" points="355" swimtime="00:04:59.48" resultid="11587" heatid="11783" lane="6" entrytime="00:05:02.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                    <SPLIT distance="100" swimtime="00:01:10.33" />
                    <SPLIT distance="150" swimtime="00:01:47.11" />
                    <SPLIT distance="200" swimtime="00:02:25.02" />
                    <SPLIT distance="250" swimtime="00:03:02.87" />
                    <SPLIT distance="300" swimtime="00:03:41.94" />
                    <SPLIT distance="350" swimtime="00:04:21.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kenzo" lastname="Kimura" birthdate="2010-04-23" gender="M" nation="BRA" license="403429" athleteid="11634" externalid="403429">
              <RESULTS>
                <RESULT eventid="1068" points="225" swimtime="00:02:43.17" resultid="11635" heatid="11724" lane="3" entrytime="00:02:43.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                    <SPLIT distance="100" swimtime="00:01:14.28" />
                    <SPLIT distance="150" swimtime="00:01:58.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="292" swimtime="00:00:30.37" resultid="11636" heatid="11764" lane="3" entrytime="00:00:32.51" entrycourse="SCM" />
                <RESULT eventid="1316" points="272" swimtime="00:01:09.13" resultid="11637" heatid="11834" lane="2" entrytime="00:01:09.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="226" swimtime="00:01:30.68" resultid="11638" heatid="11794" lane="5" entrytime="00:01:41.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Samuel" lastname="Massuda Santos" birthdate="2012-06-09" gender="M" nation="BRA" license="392189" athleteid="11626" externalid="392189">
              <RESULTS>
                <RESULT eventid="1122" points="267" swimtime="00:01:15.01" resultid="11627" heatid="11745" lane="4" entrytime="00:01:17.09" entrycourse="SCM" />
                <RESULT eventid="1170" points="299" swimtime="00:00:30.13" resultid="11628" heatid="11765" lane="1" entrytime="00:00:32.00" entrycourse="SCM" />
                <RESULT eventid="1316" points="267" swimtime="00:01:09.63" resultid="11629" heatid="11833" lane="4" entrytime="00:01:14.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1344" points="256" swimtime="00:02:52.49" resultid="11630" heatid="11848" lane="2" entrytime="00:02:59.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                    <SPLIT distance="100" swimtime="00:01:25.16" />
                    <SPLIT distance="150" swimtime="00:02:14.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Gabrieli Oliveira" birthdate="2010-09-23" gender="F" nation="BRA" license="403428" athleteid="11631" externalid="403428">
              <RESULTS>
                <RESULT eventid="1162" points="290" swimtime="00:00:34.64" resultid="11632" heatid="11760" lane="2" entrytime="00:00:33.32" entrycourse="SCM" />
                <RESULT eventid="1308" points="256" swimtime="00:01:19.09" resultid="11633" heatid="11829" lane="6" entrytime="00:01:14.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stela" lastname="Gouveia" birthdate="2014-02-27" gender="F" nation="BRA" license="415498" athleteid="11656" externalid="415498">
              <RESULTS>
                <RESULT eventid="1178" points="154" swimtime="00:00:42.73" resultid="11657" heatid="11770" lane="1" entrytime="00:00:45.22" entrycourse="SCM" />
                <RESULT eventid="1298" points="113" swimtime="00:01:43.92" resultid="11658" heatid="11820" lane="3" entrytime="00:01:56.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="117" reactiontime="+101" swimtime="00:00:51.61" resultid="11659" heatid="11800" lane="6" entrytime="00:00:51.66" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Ferreira Batista" birthdate="2014-11-26" gender="F" nation="BRA" license="392160" athleteid="11622" externalid="392160">
              <RESULTS>
                <RESULT eventid="1178" points="154" swimtime="00:00:42.75" resultid="11623" heatid="11770" lane="4" entrytime="00:00:42.40" entrycourse="SCM" />
                <RESULT eventid="1102" points="116" swimtime="00:00:58.17" resultid="11624" heatid="11735" lane="3" entrytime="00:00:58.93" entrycourse="SCM" />
                <RESULT eventid="1248" points="126" reactiontime="+51" swimtime="00:00:50.28" resultid="11625" heatid="11800" lane="2" entrytime="00:00:41.83" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Giroldo Santos" birthdate="2011-05-16" gender="M" nation="BRA" license="399602" athleteid="11639" externalid="399602">
              <RESULTS>
                <RESULT eventid="1152" points="149" swimtime="00:01:30.02" resultid="11640" heatid="11755" lane="2" entrytime="00:01:35.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="190" swimtime="00:00:35.02" resultid="11641" heatid="11764" lane="6" entrytime="00:00:34.40" entrycourse="SCM" />
                <RESULT eventid="1316" points="187" swimtime="00:01:18.28" resultid="11642" heatid="11833" lane="5" entrytime="00:01:17.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anthony" lastname="Lira Gordo" birthdate="2012-04-09" gender="M" nation="BRA" license="415261" athleteid="11652" externalid="415261">
              <RESULTS>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Tempo: 11:39)" eventid="1170" status="DSQ" swimtime="00:00:37.66" resultid="11653" heatid="11763" lane="6" entrytime="00:00:40.65" entrycourse="SCM" />
                <RESULT eventid="1316" points="134" swimtime="00:01:27.42" resultid="11654" heatid="11831" lane="3" entrytime="00:01:31.48" entrycourse="SCM" />
                <RESULT eventid="1238" points="115" swimtime="00:01:53.53" resultid="11655" heatid="11792" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique De Oliveira" birthdate="2009-07-28" gender="M" nation="BRA" license="414505" athleteid="11595" externalid="414505">
              <RESULTS>
                <RESULT eventid="1152" points="307" swimtime="00:01:10.80" resultid="11596" heatid="11756" lane="5" entrytime="00:01:13.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="363" swimtime="00:00:28.24" resultid="11597" heatid="11767" lane="6" entrytime="00:00:27.76" entrycourse="SCM" />
                <RESULT eventid="1316" points="414" swimtime="00:01:00.12" resultid="11598" heatid="11835" lane="1" entrytime="00:01:02.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rebecca" lastname="Rosa Santos" birthdate="2013-01-21" gender="F" nation="BRA" license="422158" athleteid="11675" externalid="422158">
              <RESULTS>
                <RESULT eventid="1178" points="105" swimtime="00:00:48.58" resultid="11676" heatid="11769" lane="5" entrytime="00:00:51.76" entrycourse="SCM" />
                <RESULT eventid="1298" points="77" swimtime="00:01:57.88" resultid="11677" heatid="11820" lane="6" />
                <RESULT comment="SW 6.4 - Não começou a executar a virada imediatamente após virar para a posição de peito.  (Tempo: 17:06)" eventid="1248" reactiontime="+95" status="DSQ" swimtime="00:01:03.29" resultid="11678" heatid="11798" lane="4" entrytime="00:01:05.04" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3133" nation="BRA" region="PR" clubid="11688" name="Associação Toledo Natação" shortname="Toledo Natação">
          <ATHLETES>
            <ATHLETE firstname="Arthur" lastname="Marafon Duarte" birthdate="2011-08-18" gender="M" nation="BRA" license="414184" athleteid="11689" externalid="414184">
              <RESULTS>
                <RESULT eventid="1068" points="247" swimtime="00:02:38.29" resultid="11690" heatid="11724" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                    <SPLIT distance="100" swimtime="00:01:12.14" />
                    <SPLIT distance="150" swimtime="00:01:55.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="276" swimtime="00:00:30.95" resultid="11691" heatid="11765" lane="4" entrytime="00:00:31.00" entrycourse="SCM" />
                <RESULT eventid="1316" points="253" reactiontime="+73" swimtime="00:01:10.83" resultid="11692" heatid="11834" lane="1" entrytime="00:01:10.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1214" points="167" swimtime="00:06:25.37" resultid="11693" heatid="11781" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                    <SPLIT distance="100" swimtime="00:01:29.59" />
                    <SPLIT distance="150" swimtime="00:02:18.70" />
                    <SPLIT distance="200" swimtime="00:03:07.44" />
                    <SPLIT distance="250" swimtime="00:03:56.40" />
                    <SPLIT distance="300" swimtime="00:04:45.66" />
                    <SPLIT distance="350" swimtime="00:05:36.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Torres Romancini" birthdate="2010-05-28" gender="F" nation="BRA" license="347218" athleteid="11699" externalid="347218">
              <RESULTS>
                <RESULT eventid="1112" points="409" reactiontime="+63" swimtime="00:01:13.92" resultid="11700" heatid="11742" lane="4" entrytime="00:01:13.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1162" points="436" swimtime="00:00:30.22" resultid="11701" heatid="11759" lane="6" />
                <RESULT eventid="1308" points="419" swimtime="00:01:07.12" resultid="11702" heatid="11830" lane="1" entrytime="00:01:08.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1262" points="398" reactiontime="+64" swimtime="00:02:41.60" resultid="11703" heatid="11808" lane="3" entrytime="00:02:38.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                    <SPLIT distance="100" swimtime="00:01:18.19" />
                    <SPLIT distance="150" swimtime="00:02:01.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Marafon" birthdate="2011-03-23" gender="F" nation="BRA" license="380287" athleteid="11704" externalid="380287">
              <RESULTS>
                <RESULT eventid="1086" points="354" swimtime="00:03:10.22" resultid="11705" heatid="11731" lane="1" entrytime="00:03:10.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.51" />
                    <SPLIT distance="100" swimtime="00:01:29.14" />
                    <SPLIT distance="150" swimtime="00:02:20.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1162" points="413" swimtime="00:00:30.77" resultid="11706" heatid="11761" lane="2" entrytime="00:00:30.82" entrycourse="SCM" />
                <RESULT eventid="1308" points="425" swimtime="00:01:06.83" resultid="11707" heatid="11830" lane="5" entrytime="00:01:07.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="391" swimtime="00:01:25.26" resultid="11708" heatid="11790" lane="4" entrytime="00:01:26.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Pauly Follmann" birthdate="2011-04-19" gender="F" nation="BRA" license="413886" athleteid="11709" externalid="413886">
              <RESULTS>
                <RESULT eventid="1112" points="233" reactiontime="+79" swimtime="00:01:29.08" resultid="11710" heatid="11740" lane="6" />
                <RESULT eventid="1086" points="221" swimtime="00:03:42.44" resultid="11711" heatid="11730" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.18" />
                    <SPLIT distance="100" swimtime="00:01:46.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="233" swimtime="00:01:41.31" resultid="11712" heatid="11788" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1262" points="244" reactiontime="+76" swimtime="00:03:10.16" resultid="11713" heatid="11807" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Welter Levandowski" birthdate="2011-05-06" gender="F" nation="BRA" license="380286" athleteid="11694" externalid="380286">
              <RESULTS>
                <RESULT eventid="1060" points="366" swimtime="00:02:34.15" resultid="11695" heatid="11723" lane="6" entrytime="00:02:32.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                    <SPLIT distance="100" swimtime="00:01:12.56" />
                    <SPLIT distance="150" swimtime="00:01:53.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="340" swimtime="00:11:23.39" resultid="11696" heatid="11777" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="100" swimtime="00:01:15.16" />
                    <SPLIT distance="150" swimtime="00:01:56.94" />
                    <SPLIT distance="200" swimtime="00:02:40.07" />
                    <SPLIT distance="250" swimtime="00:03:23.76" />
                    <SPLIT distance="300" swimtime="00:04:07.42" />
                    <SPLIT distance="350" swimtime="00:04:51.41" />
                    <SPLIT distance="400" swimtime="00:05:35.16" />
                    <SPLIT distance="450" swimtime="00:06:19.20" />
                    <SPLIT distance="500" swimtime="00:07:03.47" />
                    <SPLIT distance="550" swimtime="00:07:47.85" />
                    <SPLIT distance="600" swimtime="00:08:32.01" />
                    <SPLIT distance="650" swimtime="00:09:15.81" />
                    <SPLIT distance="700" swimtime="00:09:59.35" />
                    <SPLIT distance="750" swimtime="00:10:41.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="226" swimtime="00:03:16.34" resultid="11697" heatid="11812" lane="5" entrytime="00:03:19.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.26" />
                    <SPLIT distance="100" swimtime="00:01:31.53" />
                    <SPLIT distance="150" swimtime="00:02:23.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="360" swimtime="00:05:25.08" resultid="11698" heatid="11780" lane="4" entrytime="00:05:21.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                    <SPLIT distance="100" swimtime="00:01:14.43" />
                    <SPLIT distance="150" swimtime="00:01:55.39" />
                    <SPLIT distance="200" swimtime="00:02:36.95" />
                    <SPLIT distance="250" swimtime="00:03:18.95" />
                    <SPLIT distance="300" swimtime="00:04:01.39" />
                    <SPLIT distance="350" swimtime="00:04:44.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
