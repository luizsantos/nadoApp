<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.80168">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Campo Mourão" name="36º Jogos da Juventude do Paraná 2024" course="SCM" deadline="1969-12-31" hostclub="Secretaria do Esporte, Governo do Estado do Paraná" hostclub.url="https://www.esporte.pr.gov.br/" number="38325" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/newInterface/eventos/38325" startmethod="1" timing="AUTOMATIC" touchpad="ONESIDE" masters="F" state="PR" nation="BRA" hytek.courseorder="S">
      <AGEDATE value="2024-01-01" type="YEAR" />
      <POOL name="Complexo Esportivo Roberto Brzezinski" lanemin="1" lanemax="8" />
      <FACILITY city="Campo Mourão" name="Complexo Esportivo Roberto Brzezinski" nation="BRA" state="PR" street="Rua Miguel Luís Pereira" street2="Bela Vista" zip="87302-140" />
      <POINTTABLE pointtableid="3017" name="AQUA Point Scoring" version="2024" />
      <QUALIFY from="2023-01-01" until="2024-10-30" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99252-0598" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99252-0598" street="Avenida do Batel, 1230" street2="Sala 202" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2024-10-31" daytime="09:10" endtime="11:46" number="1" officialmeeting="08:30" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="1061" daytime="09:10" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2312" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1647" />
                    <RANKING order="2" place="2" resultid="1812" />
                    <RANKING order="3" place="3" resultid="1744" />
                    <RANKING order="4" place="4" resultid="1737" />
                    <RANKING order="5" place="5" resultid="1817" />
                    <RANKING order="6" place="6" resultid="1571" />
                    <RANKING order="7" place="7" resultid="1515" />
                    <RANKING order="8" place="8" resultid="1941" />
                    <RANKING order="9" place="9" resultid="1610" />
                    <RANKING order="10" place="10" resultid="2056" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2358" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2359" daytime="09:34" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1074" daytime="10:00" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2313" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1519" />
                    <RANKING order="2" place="2" resultid="1539" />
                    <RANKING order="3" place="3" resultid="1642" />
                    <RANKING order="4" place="4" resultid="1634" />
                    <RANKING order="5" place="5" resultid="1911" />
                    <RANKING order="6" place="6" resultid="1560" />
                    <RANKING order="7" place="7" resultid="1871" />
                    <RANKING order="8" place="8" resultid="1765" />
                    <RANKING order="9" place="9" resultid="1787" />
                    <RANKING order="10" place="10" resultid="2045" />
                    <RANKING order="11" place="11" resultid="1778" />
                    <RANKING order="12" place="12" resultid="1938" />
                    <RANKING order="13" place="-1" resultid="1704" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2360" daytime="10:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2361" daytime="10:04" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1087" daytime="10:08" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2314" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1555" />
                    <RANKING order="2" place="2" resultid="1529" />
                    <RANKING order="3" place="3" resultid="1755" />
                    <RANKING order="4" place="4" resultid="1593" />
                    <RANKING order="5" place="5" resultid="1896" />
                    <RANKING order="6" place="6" resultid="1714" />
                    <RANKING order="7" place="7" resultid="1701" />
                    <RANKING order="8" place="8" resultid="2022" />
                    <RANKING order="9" place="9" resultid="1963" />
                    <RANKING order="10" place="10" resultid="1931" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2362" daytime="10:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2363" daytime="10:12" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1100" daytime="10:18" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2316" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1672" />
                    <RANKING order="2" place="2" resultid="1643" />
                    <RANKING order="3" place="3" resultid="1844" />
                    <RANKING order="4" place="4" resultid="1579" />
                    <RANKING order="5" place="5" resultid="1876" />
                    <RANKING order="6" place="6" resultid="1861" />
                    <RANKING order="7" place="7" resultid="1598" />
                    <RANKING order="8" place="8" resultid="1924" />
                    <RANKING order="9" place="9" resultid="2025" />
                    <RANKING order="10" place="10" resultid="2065" />
                    <RANKING order="11" place="11" resultid="1807" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2364" daytime="10:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2365" daytime="10:20" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1113" daytime="10:22" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2318" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1638" />
                    <RANKING order="2" place="2" resultid="1995" />
                    <RANKING order="3" place="3" resultid="1530" />
                    <RANKING order="4" place="4" resultid="2050" />
                    <RANKING order="5" place="5" resultid="1952" />
                    <RANKING order="6" place="6" resultid="1731" />
                    <RANKING order="7" place="7" resultid="1901" />
                    <RANKING order="8" place="8" resultid="1719" />
                    <RANKING order="9" place="8" resultid="1825" />
                    <RANKING order="10" place="10" resultid="1783" />
                    <RANKING order="11" place="11" resultid="2070" />
                    <RANKING order="12" place="-1" resultid="1940" />
                    <RANKING order="13" place="-1" resultid="2000" />
                    <RANKING order="14" place="-1" resultid="2003" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2366" daytime="10:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2367" daytime="10:26" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1126" daytime="10:42" gender="M" number="6" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2317" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1865" />
                    <RANKING order="2" place="2" resultid="2350" />
                    <RANKING order="3" place="3" resultid="1657" />
                    <RANKING order="4" place="3" resultid="1984" />
                    <RANKING order="5" place="5" resultid="1689" />
                    <RANKING order="6" place="6" resultid="2012" />
                    <RANKING order="7" place="7" resultid="1875" />
                    <RANKING order="8" place="8" resultid="1860" />
                    <RANKING order="9" place="9" resultid="1497" />
                    <RANKING order="10" place="10" resultid="1764" />
                    <RANKING order="11" place="10" resultid="1834" />
                    <RANKING order="12" place="12" resultid="2017" />
                    <RANKING order="13" place="13" resultid="1849" />
                    <RANKING order="14" place="14" resultid="1543" />
                    <RANKING order="15" place="15" resultid="2044" />
                    <RANKING order="16" place="16" resultid="1606" />
                    <RANKING order="17" place="17" resultid="1489" />
                    <RANKING order="18" place="18" resultid="1575" />
                    <RANKING order="19" place="19" resultid="1505" />
                    <RANKING order="20" place="20" resultid="2079" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2368" daytime="10:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2369" daytime="10:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2370" daytime="10:46" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1139" daytime="10:50" gender="F" number="7" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2320" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1652" />
                    <RANKING order="2" place="2" resultid="1709" />
                    <RANKING order="3" place="3" resultid="1994" />
                    <RANKING order="4" place="4" resultid="1743" />
                    <RANKING order="5" place="5" resultid="1821" />
                    <RANKING order="6" place="6" resultid="1619" />
                    <RANKING order="7" place="7" resultid="1782" />
                    <RANKING order="8" place="8" resultid="1534" />
                    <RANKING order="9" place="9" resultid="1906" />
                    <RANKING order="10" place="10" resultid="1570" />
                    <RANKING order="11" place="11" resultid="1920" />
                    <RANKING order="12" place="12" resultid="1934" />
                    <RANKING order="13" place="13" resultid="1502" />
                    <RANKING order="14" place="14" resultid="2034" />
                    <RANKING order="15" place="15" resultid="1802" />
                    <RANKING order="16" place="-1" resultid="1999" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2371" daytime="10:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2372" daytime="10:52" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1152" daytime="10:54" gender="M" number="8" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2322" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1524" />
                    <RANKING order="2" place="2" resultid="1602" />
                    <RANKING order="3" place="3" resultid="1667" />
                    <RANKING order="4" place="4" resultid="1551" />
                    <RANKING order="5" place="5" resultid="1633" />
                    <RANKING order="6" place="6" resultid="1681" />
                    <RANKING order="7" place="7" resultid="1916" />
                    <RANKING order="8" place="8" resultid="1989" />
                    <RANKING order="9" place="9" resultid="1870" />
                    <RANKING order="10" place="10" resultid="1829" />
                    <RANKING order="11" place="11" resultid="1792" />
                    <RANKING order="12" place="12" resultid="1777" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2373" daytime="10:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2374" daytime="10:58" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1165" daytime="11:04" gender="F" number="9" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2321" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1759" />
                    <RANKING order="2" place="2" resultid="1653" />
                    <RANKING order="3" place="3" resultid="1565" />
                    <RANKING order="4" place="4" resultid="1754" />
                    <RANKING order="5" place="5" resultid="1514" />
                    <RANKING order="6" place="6" resultid="1692" />
                    <RANKING order="7" place="7" resultid="1945" />
                    <RANKING order="8" place="8" resultid="1588" />
                    <RANKING order="9" place="9" resultid="2055" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2375" daytime="11:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2376" daytime="11:08" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1178" daytime="11:14" gender="M" number="10" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2323" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2351" />
                    <RANKING order="2" place="2" resultid="1912" />
                    <RANKING order="3" place="3" resultid="1727" />
                    <RANKING order="4" place="4" resultid="1705" />
                    <RANKING order="5" place="5" resultid="1547" />
                    <RANKING order="6" place="6" resultid="1928" />
                    <RANKING order="7" place="7" resultid="1880" />
                    <RANKING order="8" place="8" resultid="2026" />
                    <RANKING order="9" place="9" resultid="1561" />
                    <RANKING order="10" place="10" resultid="1498" />
                    <RANKING order="11" place="11" resultid="1615" />
                    <RANKING order="12" place="12" resultid="1850" />
                    <RANKING order="13" place="13" resultid="2075" />
                    <RANKING order="14" place="14" resultid="1808" />
                    <RANKING order="15" place="15" resultid="1494" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2377" daytime="11:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2378" daytime="11:16" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1191" daytime="11:18" gender="F" number="11" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2324" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1978" />
                    <RANKING order="2" place="2" resultid="1897" />
                    <RANKING order="3" place="3" resultid="1696" />
                    <RANKING order="4" place="4" resultid="2060" />
                    <RANKING order="5" place="5" resultid="2008" />
                    <RANKING order="6" place="6" resultid="1892" />
                    <RANKING order="7" place="7" resultid="1715" />
                    <RANKING order="8" place="8" resultid="1594" />
                    <RANKING order="9" place="9" resultid="1822" />
                    <RANKING order="10" place="10" resultid="1589" />
                    <RANKING order="11" place="11" resultid="1964" />
                    <RANKING order="12" place="12" resultid="2030" />
                    <RANKING order="13" place="13" resultid="2071" />
                    <RANKING order="14" place="-1" resultid="1803" />
                    <RANKING order="15" place="-1" resultid="2035" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2379" daytime="11:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2380" daytime="11:20" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1204" daytime="11:38" gender="X" number="12" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1205" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1857" />
                    <RANKING order="2" place="2" resultid="1627" />
                    <RANKING order="3" place="3" resultid="2085" />
                    <RANKING order="4" place="-1" resultid="1751" />
                    <RANKING order="5" place="-1" resultid="1974" />
                    <RANKING order="6" place="-1" resultid="2041" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2381" daytime="11:38" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-10-31" daytime="16:10" endtime="19:15" number="2" officialmeeting="15:30" warmupfrom="15:00" warmupuntil="16:00">
          <EVENTS>
            <EVENT eventid="1206" daytime="16:10" gender="F" number="13" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2325" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1760" />
                    <RANKING order="2" place="2" resultid="1648" />
                    <RANKING order="3" place="3" resultid="1566" />
                    <RANKING order="4" place="4" resultid="1693" />
                    <RANKING order="5" place="5" resultid="1738" />
                    <RANKING order="6" place="6" resultid="1814" />
                    <RANKING order="7" place="7" resultid="1612" />
                    <RANKING order="8" place="8" resultid="1946" />
                    <RANKING order="9" place="9" resultid="1818" />
                    <RANKING order="10" place="10" resultid="1572" />
                    <RANKING order="11" place="11" resultid="2058" />
                    <RANKING order="12" place="12" resultid="1903" />
                    <RANKING order="13" place="13" resultid="1935" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2382" daytime="16:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2383" daytime="16:18" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1219" daytime="16:24" gender="M" number="14" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2326" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1520" />
                    <RANKING order="2" place="2" resultid="1658" />
                    <RANKING order="3" place="3" resultid="1525" />
                    <RANKING order="4" place="4" resultid="1985" />
                    <RANKING order="5" place="5" resultid="1867" />
                    <RANKING order="6" place="6" resultid="1723" />
                    <RANKING order="7" place="7" resultid="1544" />
                    <RANKING order="8" place="8" resultid="1793" />
                    <RANKING order="9" place="9" resultid="2018" />
                    <RANKING order="10" place="10" resultid="1885" />
                    <RANKING order="11" place="11" resultid="1789" />
                    <RANKING order="12" place="12" resultid="1968" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2384" daytime="16:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2385" daytime="16:30" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1232" daytime="16:38" gender="F" number="15" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2327" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1595" />
                    <RANKING order="2" place="2" resultid="1556" />
                    <RANKING order="3" place="3" resultid="1979" />
                    <RANKING order="4" place="4" resultid="1697" />
                    <RANKING order="5" place="5" resultid="1898" />
                    <RANKING order="6" place="6" resultid="1716" />
                    <RANKING order="7" place="7" resultid="1590" />
                    <RANKING order="8" place="8" resultid="2061" />
                    <RANKING order="9" place="9" resultid="2009" />
                    <RANKING order="10" place="10" resultid="1840" />
                    <RANKING order="11" place="11" resultid="1965" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2386" daytime="16:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2387" daytime="16:42" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1245" daytime="16:48" gender="M" number="16" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2328" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1990" />
                    <RANKING order="2" place="2" resultid="1913" />
                    <RANKING order="3" place="3" resultid="1728" />
                    <RANKING order="4" place="4" resultid="1630" />
                    <RANKING order="5" place="5" resultid="1772" />
                    <RANKING order="6" place="6" resultid="1583" />
                    <RANKING order="7" place="7" resultid="1706" />
                    <RANKING order="8" place="8" resultid="1881" />
                    <RANKING order="9" place="9" resultid="1616" />
                    <RANKING order="10" place="10" resultid="1576" />
                    <RANKING order="11" place="11" resultid="1797" />
                    <RANKING order="12" place="12" resultid="1890" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2388" daytime="16:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2389" daytime="16:52" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1258" daytime="16:56" gender="F" number="17" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2331" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1655" />
                    <RANKING order="2" place="2" resultid="1711" />
                    <RANKING order="3" place="3" resultid="1823" />
                    <RANKING order="4" place="4" resultid="1954" />
                    <RANKING order="5" place="5" resultid="1784" />
                    <RANKING order="6" place="6" resultid="1893" />
                    <RANKING order="7" place="7" resultid="2062" />
                    <RANKING order="8" place="8" resultid="1620" />
                    <RANKING order="9" place="9" resultid="1908" />
                    <RANKING order="10" place="10" resultid="2036" />
                    <RANKING order="11" place="11" resultid="1804" />
                    <RANKING order="12" place="12" resultid="1503" />
                    <RANKING order="13" place="-1" resultid="2072" />
                    <RANKING order="14" place="-1" resultid="2001" />
                    <RANKING order="15" place="-1" resultid="2005" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2390" daytime="16:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2391" daytime="16:58" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1271" daytime="17:00" gender="M" number="18" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2329" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1665" />
                    <RANKING order="2" place="2" resultid="1659" />
                    <RANKING order="3" place="3" resultid="1986" />
                    <RANKING order="4" place="4" resultid="1877" />
                    <RANKING order="5" place="5" resultid="1678" />
                    <RANKING order="6" place="6" resultid="1766" />
                    <RANKING order="7" place="7" resultid="2014" />
                    <RANKING order="8" place="8" resultid="1863" />
                    <RANKING order="9" place="9" resultid="1499" />
                    <RANKING order="10" place="10" resultid="1562" />
                    <RANKING order="11" place="11" resultid="2046" />
                    <RANKING order="12" place="12" resultid="1851" />
                    <RANKING order="13" place="13" resultid="1846" />
                    <RANKING order="14" place="14" resultid="2027" />
                    <RANKING order="15" place="15" resultid="1491" />
                    <RANKING order="16" place="16" resultid="1957" />
                    <RANKING order="17" place="17" resultid="2081" />
                    <RANKING order="18" place="18" resultid="1506" />
                    <RANKING order="19" place="-1" resultid="1584" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2392" daytime="17:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2393" daytime="17:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2394" daytime="17:04" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1284" daytime="17:20" gender="F" number="19" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2330" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1639" />
                    <RANKING order="2" place="2" resultid="1531" />
                    <RANKING order="3" place="3" resultid="1996" />
                    <RANKING order="4" place="4" resultid="1535" />
                    <RANKING order="5" place="5" resultid="2051" />
                    <RANKING order="6" place="6" resultid="1732" />
                    <RANKING order="7" place="7" resultid="1720" />
                    <RANKING order="8" place="8" resultid="1942" />
                    <RANKING order="9" place="9" resultid="1611" />
                    <RANKING order="10" place="10" resultid="1826" />
                    <RANKING order="11" place="11" resultid="1902" />
                    <RANKING order="12" place="12" resultid="1813" />
                    <RANKING order="13" place="13" resultid="1839" />
                    <RANKING order="14" place="-1" resultid="2004" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2395" daytime="17:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2396" daytime="17:26" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1297" daytime="17:30" gender="M" number="20" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2333" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1673" />
                    <RANKING order="2" place="2" resultid="1540" />
                    <RANKING order="3" place="3" resultid="1835" />
                    <RANKING order="4" place="4" resultid="1685" />
                    <RANKING order="5" place="5" resultid="1662" />
                    <RANKING order="6" place="6" resultid="1599" />
                    <RANKING order="7" place="7" resultid="1845" />
                    <RANKING order="8" place="8" resultid="1925" />
                    <RANKING order="9" place="9" resultid="1862" />
                    <RANKING order="10" place="10" resultid="1788" />
                    <RANKING order="11" place="11" resultid="1607" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2397" daytime="17:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2398" daytime="17:36" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1310" daytime="17:40" gender="F" number="21" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2335" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1654" />
                    <RANKING order="2" place="2" resultid="1756" />
                    <RANKING order="3" place="3" resultid="1710" />
                    <RANKING order="4" place="4" resultid="1745" />
                    <RANKING order="5" place="5" resultid="1516" />
                    <RANKING order="6" place="6" resultid="1769" />
                    <RANKING order="7" place="7" resultid="1907" />
                    <RANKING order="8" place="8" resultid="2057" />
                    <RANKING order="9" place="-1" resultid="1953" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2399" daytime="17:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2400" daytime="17:42" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1323" daytime="17:46" gender="M" number="22" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2336" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1866" />
                    <RANKING order="2" place="2" resultid="1872" />
                    <RANKING order="3" place="3" resultid="1603" />
                    <RANKING order="4" place="4" resultid="1644" />
                    <RANKING order="5" place="5" resultid="1580" />
                    <RANKING order="6" place="6" resultid="2013" />
                    <RANKING order="7" place="7" resultid="1682" />
                    <RANKING order="8" place="8" resultid="1917" />
                    <RANKING order="9" place="9" resultid="1668" />
                    <RANKING order="10" place="10" resultid="1552" />
                    <RANKING order="11" place="11" resultid="1830" />
                    <RANKING order="12" place="12" resultid="1779" />
                    <RANKING order="13" place="13" resultid="1490" />
                    <RANKING order="14" place="14" resultid="1809" />
                    <RANKING order="15" place="15" resultid="1508" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2401" daytime="17:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2402" daytime="17:48" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1336" daytime="17:52" gender="F" number="23" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2338" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1761" />
                    <RANKING order="2" place="2" resultid="1557" />
                    <RANKING order="3" place="3" resultid="1649" />
                    <RANKING order="4" place="4" resultid="1567" />
                    <RANKING order="5" place="5" resultid="1536" />
                    <RANKING order="6" place="6" resultid="1980" />
                    <RANKING order="7" place="7" resultid="1702" />
                    <RANKING order="8" place="8" resultid="1947" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2403" daytime="17:52" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1349" daytime="18:00" gender="M" number="24" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2340" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1521" />
                    <RANKING order="2" place="2" resultid="1526" />
                    <RANKING order="3" place="3" resultid="1773" />
                    <RANKING order="4" place="4" resultid="1548" />
                    <RANKING order="5" place="5" resultid="1724" />
                    <RANKING order="6" place="6" resultid="1991" />
                    <RANKING order="7" place="7" resultid="1635" />
                    <RANKING order="8" place="8" resultid="1740" />
                    <RANKING order="9" place="9" resultid="1882" />
                    <RANKING order="10" place="10" resultid="1799" />
                    <RANKING order="11" place="-1" resultid="1886" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2404" daytime="18:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2405" daytime="18:08" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1362" daytime="18:30" gender="F" number="25" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1363" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1747" />
                    <RANKING order="2" place="2" resultid="1853" />
                    <RANKING order="3" place="3" resultid="1623" />
                    <RANKING order="4" place="4" resultid="1970" />
                    <RANKING order="5" place="5" resultid="2037" />
                    <RANKING order="6" place="6" resultid="2083" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2406" daytime="18:30" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1364" daytime="18:38" gender="M" number="26" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1365" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1749" />
                    <RANKING order="2" place="2" resultid="1972" />
                    <RANKING order="3" place="3" resultid="1625" />
                    <RANKING order="4" place="4" resultid="1855" />
                    <RANKING order="5" place="5" resultid="2039" />
                    <RANKING order="6" place="6" resultid="1510" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2407" daytime="18:38" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-11-01" daytime="09:10" endtime="11:25" number="3" officialmeeting="08:30" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="1366" daytime="09:10" gender="F" number="27" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2341" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1640" />
                    <RANKING order="2" place="2" resultid="1532" />
                    <RANKING order="3" place="3" resultid="2052" />
                    <RANKING order="4" place="4" resultid="1997" />
                    <RANKING order="5" place="5" resultid="1733" />
                    <RANKING order="6" place="6" resultid="1943" />
                    <RANKING order="7" place="7" resultid="1537" />
                    <RANKING order="8" place="8" resultid="1955" />
                    <RANKING order="9" place="9" resultid="1721" />
                    <RANKING order="10" place="10" resultid="1904" />
                    <RANKING order="11" place="11" resultid="1827" />
                    <RANKING order="12" place="12" resultid="1841" />
                    <RANKING order="13" place="13" resultid="1621" />
                    <RANKING order="14" place="14" resultid="1785" />
                    <RANKING order="15" place="15" resultid="2023" />
                    <RANKING order="16" place="-1" resultid="2006" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2408" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2409" daytime="09:14" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1379" daytime="09:16" gender="M" number="28" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2343" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1645" />
                    <RANKING order="2" place="2" resultid="1636" />
                    <RANKING order="3" place="3" resultid="1581" />
                    <RANKING order="4" place="4" resultid="1836" />
                    <RANKING order="5" place="5" resultid="1847" />
                    <RANKING order="6" place="6" resultid="1600" />
                    <RANKING order="7" place="7" resultid="1878" />
                    <RANKING order="8" place="8" resultid="1926" />
                    <RANKING order="9" place="9" resultid="1790" />
                    <RANKING order="10" place="10" resultid="1608" />
                    <RANKING order="11" place="11" resultid="1950" />
                    <RANKING order="12" place="-1" resultid="1674" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2410" daytime="09:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2411" daytime="09:20" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1392" daytime="09:24" gender="F" number="29" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2342" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1762" />
                    <RANKING order="2" place="2" resultid="1650" />
                    <RANKING order="3" place="3" resultid="1746" />
                    <RANKING order="4" place="4" resultid="1613" />
                    <RANKING order="5" place="5" resultid="1815" />
                    <RANKING order="6" place="6" resultid="1819" />
                    <RANKING order="7" place="7" resultid="1573" />
                    <RANKING order="8" place="8" resultid="1622" />
                    <RANKING order="9" place="9" resultid="1676" />
                    <RANKING order="10" place="10" resultid="1936" />
                    <RANKING order="11" place="11" resultid="1932" />
                    <RANKING order="12" place="12" resultid="1921" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2412" daytime="09:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2413" daytime="09:28" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1405" daytime="09:32" gender="M" number="30" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2344" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1987" />
                    <RANKING order="2" place="2" resultid="1660" />
                    <RANKING order="3" place="3" resultid="1775" />
                    <RANKING order="4" place="4" resultid="1687" />
                    <RANKING order="5" place="5" resultid="1586" />
                    <RANKING order="6" place="6" resultid="1690" />
                    <RANKING order="7" place="7" resultid="1553" />
                    <RANKING order="8" place="8" resultid="2020" />
                    <RANKING order="9" place="9" resultid="1888" />
                    <RANKING order="10" place="10" resultid="2047" />
                    <RANKING order="11" place="11" resultid="1958" />
                    <RANKING order="12" place="12" resultid="1563" />
                    <RANKING order="13" place="13" resultid="1795" />
                    <RANKING order="14" place="14" resultid="1831" />
                    <RANKING order="15" place="-1" resultid="1868" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2414" daytime="09:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2415" daytime="09:36" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1418" daytime="09:40" gender="F" number="31" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2345" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1757" />
                    <RANKING order="2" place="2" resultid="1712" />
                    <RANKING order="3" place="3" resultid="1770" />
                    <RANKING order="4" place="4" resultid="1948" />
                    <RANKING order="5" place="5" resultid="1517" />
                    <RANKING order="6" place="6" resultid="1909" />
                    <RANKING order="7" place="7" resultid="1568" />
                    <RANKING order="8" place="8" resultid="1694" />
                    <RANKING order="9" place="9" resultid="2053" />
                    <RANKING order="10" place="10" resultid="1922" />
                    <RANKING order="11" place="11" resultid="1805" />
                    <RANKING order="12" place="-1" resultid="1735" />
                    <RANKING order="13" place="-1" resultid="2032" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2416" daytime="09:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2417" daytime="09:42" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1431" daytime="09:44" gender="M" number="32" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2346" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1873" />
                    <RANKING order="2" place="2" resultid="1679" />
                    <RANKING order="3" place="3" resultid="1683" />
                    <RANKING order="4" place="4" resultid="1918" />
                    <RANKING order="5" place="5" resultid="2015" />
                    <RANKING order="6" place="6" resultid="1670" />
                    <RANKING order="7" place="7" resultid="1604" />
                    <RANKING order="8" place="8" resultid="1767" />
                    <RANKING order="9" place="9" resultid="1492" />
                    <RANKING order="10" place="10" resultid="1959" />
                    <RANKING order="11" place="11" resultid="1837" />
                    <RANKING order="12" place="12" resultid="1832" />
                    <RANKING order="13" place="13" resultid="1545" />
                    <RANKING order="14" place="14" resultid="1577" />
                    <RANKING order="15" place="15" resultid="1509" />
                    <RANKING order="16" place="16" resultid="2082" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2418" daytime="09:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2419" daytime="09:46" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1444" daytime="10:02" gender="F" number="33" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2347" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1981" />
                    <RANKING order="2" place="2" resultid="1899" />
                    <RANKING order="3" place="3" resultid="1558" />
                    <RANKING order="4" place="4" resultid="1698" />
                    <RANKING order="5" place="5" resultid="2010" />
                    <RANKING order="6" place="6" resultid="1717" />
                    <RANKING order="7" place="7" resultid="1596" />
                    <RANKING order="8" place="8" resultid="2429" />
                    <RANKING order="9" place="9" resultid="1591" />
                    <RANKING order="10" place="10" resultid="1842" />
                    <RANKING order="11" place="11" resultid="1894" />
                    <RANKING order="12" place="12" resultid="1966" />
                    <RANKING order="13" place="13" resultid="2031" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2420" daytime="10:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2421" daytime="10:06" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1457" daytime="10:08" gender="M" number="34" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2348" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1729" />
                    <RANKING order="2" place="2" resultid="1914" />
                    <RANKING order="3" place="3" resultid="1992" />
                    <RANKING order="4" place="4" resultid="1707" />
                    <RANKING order="5" place="5" resultid="1549" />
                    <RANKING order="6" place="6" resultid="1631" />
                    <RANKING order="7" place="7" resultid="1883" />
                    <RANKING order="8" place="8" resultid="1929" />
                    <RANKING order="9" place="9" resultid="1617" />
                    <RANKING order="10" place="10" resultid="1500" />
                    <RANKING order="11" place="11" resultid="2028" />
                    <RANKING order="12" place="12" resultid="1585" />
                    <RANKING order="13" place="13" resultid="1800" />
                    <RANKING order="14" place="14" resultid="1852" />
                    <RANKING order="15" place="15" resultid="2077" />
                    <RANKING order="16" place="16" resultid="1495" />
                    <RANKING order="17" place="-1" resultid="1810" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2422" daytime="10:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2423" daytime="10:12" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2424" daytime="10:14" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1470" daytime="10:16" gender="M" number="35" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2349" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1522" />
                    <RANKING order="2" place="2" resultid="1527" />
                    <RANKING order="3" place="3" resultid="1774" />
                    <RANKING order="4" place="4" resultid="1725" />
                    <RANKING order="5" place="5" resultid="1541" />
                    <RANKING order="6" place="6" resultid="1686" />
                    <RANKING order="7" place="7" resultid="1741" />
                    <RANKING order="8" place="8" resultid="1887" />
                    <RANKING order="9" place="9" resultid="2019" />
                    <RANKING order="10" place="10" resultid="1780" />
                    <RANKING order="11" place="11" resultid="1969" />
                    <RANKING order="12" place="12" resultid="1794" />
                    <RANKING order="13" place="13" resultid="1961" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2425" daytime="10:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2426" daytime="10:30" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1483" daytime="10:56" gender="F" number="36" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1484" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1748" />
                    <RANKING order="2" place="2" resultid="1624" />
                    <RANKING order="3" place="3" resultid="1854" />
                    <RANKING order="4" place="4" resultid="1971" />
                    <RANKING order="5" place="5" resultid="2038" />
                    <RANKING order="6" place="-1" resultid="2084" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2427" daytime="10:56" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1485" daytime="11:04" gender="M" number="37" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1486" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1973" />
                    <RANKING order="2" place="2" resultid="1626" />
                    <RANKING order="3" place="3" resultid="1511" />
                    <RANKING order="4" place="-1" resultid="1750" />
                    <RANKING order="5" place="-1" resultid="2040" />
                    <RANKING order="6" place="-1" resultid="1856" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2428" daytime="11:04" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="1492" nation="BRA" region="PR" clubid="1628" name="Seleção De Curitiba/PR" shortname="Curitiba">
          <ATHLETES>
            <ATHLETE firstname="Julia" lastname="Nalle Bejes" birthdate="2010-04-20" gender="F" nation="BRA" license="377323" athleteid="1700" externalid="377323">
              <RESULTS>
                <RESULT eventid="1087" points="330" swimtime="00:02:56.22" resultid="1701" heatid="2362" lane="5" entrytime="00:03:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.85" />
                    <SPLIT distance="100" swimtime="00:01:27.41" />
                    <SPLIT distance="150" swimtime="00:02:15.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="340" swimtime="00:06:10.72" resultid="1702" heatid="2403" lane="1" entrytime="00:06:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.13" />
                    <SPLIT distance="100" swimtime="00:01:31.39" />
                    <SPLIT distance="150" swimtime="00:02:20.06" />
                    <SPLIT distance="200" swimtime="00:03:09.00" />
                    <SPLIT distance="250" swimtime="00:03:55.80" />
                    <SPLIT distance="300" swimtime="00:04:45.94" />
                    <SPLIT distance="350" swimtime="00:05:30.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lauren" lastname="Dziura" birthdate="2010-01-11" gender="F" nation="BRA" license="369416" athleteid="1736" externalid="369416">
              <RESULTS>
                <RESULT eventid="1061" points="419" swimtime="00:20:13.41" resultid="1737" heatid="2358" lane="3" entrytime="00:23:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.57" />
                    <SPLIT distance="300" swimtime="00:03:51.20" />
                    <SPLIT distance="350" swimtime="00:04:31.56" />
                    <SPLIT distance="400" swimtime="00:05:11.73" />
                    <SPLIT distance="450" swimtime="00:05:52.10" />
                    <SPLIT distance="500" swimtime="00:06:32.91" />
                    <SPLIT distance="550" swimtime="00:07:13.65" />
                    <SPLIT distance="600" swimtime="00:07:54.87" />
                    <SPLIT distance="650" swimtime="00:08:35.40" />
                    <SPLIT distance="700" swimtime="00:09:16.57" />
                    <SPLIT distance="750" swimtime="00:09:57.64" />
                    <SPLIT distance="800" swimtime="00:10:38.36" />
                    <SPLIT distance="850" swimtime="00:11:20.15" />
                    <SPLIT distance="900" swimtime="00:12:00.92" />
                    <SPLIT distance="950" swimtime="00:12:42.75" />
                    <SPLIT distance="1000" swimtime="00:13:23.92" />
                    <SPLIT distance="1050" swimtime="00:14:04.92" />
                    <SPLIT distance="1100" swimtime="00:14:46.23" />
                    <SPLIT distance="1150" swimtime="00:15:27.23" />
                    <SPLIT distance="1200" swimtime="00:16:09.52" />
                    <SPLIT distance="1250" swimtime="00:16:51.17" />
                    <SPLIT distance="1300" swimtime="00:17:31.97" />
                    <SPLIT distance="1350" swimtime="00:18:13.07" />
                    <SPLIT distance="1400" swimtime="00:18:53.58" />
                    <SPLIT distance="1450" swimtime="00:20:13.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="450" swimtime="00:05:01.69" resultid="1738" heatid="2382" lane="5" entrytime="00:05:12.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                    <SPLIT distance="100" swimtime="00:01:12.78" />
                    <SPLIT distance="150" swimtime="00:01:50.79" />
                    <SPLIT distance="200" swimtime="00:02:29.31" />
                    <SPLIT distance="250" swimtime="00:03:07.77" />
                    <SPLIT distance="300" swimtime="00:03:45.87" />
                    <SPLIT distance="350" swimtime="00:04:24.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabelly" lastname="Sinnott" birthdate="2009-03-14" gender="F" nation="BRA" license="367255" athleteid="1646" externalid="367255">
              <RESULTS>
                <RESULT eventid="1061" points="562" swimtime="00:18:20.51" resultid="1647" heatid="2359" lane="4" entrytime="00:18:34.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="100" swimtime="00:01:09.37" />
                    <SPLIT distance="150" swimtime="00:01:45.49" />
                    <SPLIT distance="200" swimtime="00:02:22.02" />
                    <SPLIT distance="250" swimtime="00:02:58.77" />
                    <SPLIT distance="300" swimtime="00:03:35.38" />
                    <SPLIT distance="350" swimtime="00:04:12.12" />
                    <SPLIT distance="400" swimtime="00:04:48.75" />
                    <SPLIT distance="450" swimtime="00:05:25.63" />
                    <SPLIT distance="500" swimtime="00:06:02.37" />
                    <SPLIT distance="550" swimtime="00:06:39.25" />
                    <SPLIT distance="600" swimtime="00:07:16.23" />
                    <SPLIT distance="650" swimtime="00:07:52.73" />
                    <SPLIT distance="700" swimtime="00:08:29.96" />
                    <SPLIT distance="750" swimtime="00:09:07.07" />
                    <SPLIT distance="800" swimtime="00:09:43.71" />
                    <SPLIT distance="850" swimtime="00:10:20.61" />
                    <SPLIT distance="900" swimtime="00:10:57.82" />
                    <SPLIT distance="950" swimtime="00:11:34.93" />
                    <SPLIT distance="1000" swimtime="00:12:11.83" />
                    <SPLIT distance="1050" swimtime="00:12:48.75" />
                    <SPLIT distance="1100" swimtime="00:13:25.70" />
                    <SPLIT distance="1150" swimtime="00:14:03.13" />
                    <SPLIT distance="1200" swimtime="00:14:40.00" />
                    <SPLIT distance="1250" swimtime="00:15:17.27" />
                    <SPLIT distance="1300" swimtime="00:15:54.11" />
                    <SPLIT distance="1350" swimtime="00:16:31.26" />
                    <SPLIT distance="1400" swimtime="00:17:08.89" />
                    <SPLIT distance="1450" swimtime="00:17:45.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="583" swimtime="00:04:36.73" resultid="1648" heatid="2383" lane="4" entrytime="00:04:40.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                    <SPLIT distance="100" swimtime="00:01:05.98" />
                    <SPLIT distance="150" swimtime="00:01:40.40" />
                    <SPLIT distance="200" swimtime="00:02:15.34" />
                    <SPLIT distance="250" swimtime="00:02:50.65" />
                    <SPLIT distance="300" swimtime="00:03:26.19" />
                    <SPLIT distance="350" swimtime="00:04:01.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="465" swimtime="00:05:34.19" resultid="1649" heatid="2403" lane="3" entrytime="00:05:41.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                    <SPLIT distance="100" swimtime="00:01:14.32" />
                    <SPLIT distance="150" swimtime="00:01:59.98" />
                    <SPLIT distance="200" swimtime="00:02:42.95" />
                    <SPLIT distance="250" swimtime="00:03:31.89" />
                    <SPLIT distance="300" swimtime="00:04:21.46" />
                    <SPLIT distance="350" swimtime="00:04:58.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="608" swimtime="00:02:10.18" resultid="1650" heatid="2412" lane="5" entrytime="00:02:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                    <SPLIT distance="100" swimtime="00:01:02.87" />
                    <SPLIT distance="150" swimtime="00:01:36.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabelly" lastname="Mendonca Bello" birthdate="2008-04-15" gender="F" nation="BRA" license="376996" athleteid="1713" externalid="376996" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1087" points="398" swimtime="00:02:45.66" resultid="1714" heatid="2363" lane="7" entrytime="00:02:55.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                    <SPLIT distance="100" swimtime="00:01:20.78" />
                    <SPLIT distance="150" swimtime="00:02:07.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="390" swimtime="00:00:38.83" resultid="1715" heatid="2380" lane="1" entrytime="00:00:40.84" entrycourse="SCM" />
                <RESULT eventid="1232" points="430" swimtime="00:02:58.17" resultid="1716" heatid="2387" lane="2" entrytime="00:03:10.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.89" />
                    <SPLIT distance="100" swimtime="00:01:26.44" />
                    <SPLIT distance="150" swimtime="00:02:12.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1444" points="405" swimtime="00:01:24.23" resultid="1717" heatid="2421" lane="6" entrytime="00:01:24.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ricardo" lastname="De Lima Cavalcanti" birthdate="2009-12-17" gender="M" nation="BRA" license="380965" athleteid="1666" externalid="380965">
              <RESULTS>
                <RESULT eventid="1152" points="432" swimtime="00:02:21.34" resultid="1667" heatid="2374" lane="3" entrytime="00:02:22.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                    <SPLIT distance="100" swimtime="00:01:06.55" />
                    <SPLIT distance="150" swimtime="00:01:44.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1323" points="391" swimtime="00:01:05.32" resultid="1668" heatid="2402" lane="6" entrytime="00:01:01.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" status="RJC" swimtime="00:00:00.00" resultid="1669" />
                <RESULT eventid="1431" points="429" swimtime="00:00:28.83" resultid="1670" heatid="2419" lane="7" entrytime="00:00:28.60" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jhon" lastname="Caleb Dos Santos" birthdate="2010-03-02" gender="M" nation="BRA" license="359020" athleteid="1632" externalid="359020">
              <RESULTS>
                <RESULT eventid="1152" points="421" swimtime="00:02:22.48" resultid="1633" heatid="2373" lane="5" entrytime="00:03:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                    <SPLIT distance="100" swimtime="00:01:08.11" />
                    <SPLIT distance="150" swimtime="00:01:45.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="473" swimtime="00:02:20.69" resultid="1634" heatid="2361" lane="6" entrytime="00:02:20.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.33" />
                    <SPLIT distance="100" swimtime="00:01:06.23" />
                    <SPLIT distance="150" swimtime="00:01:47.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="415" swimtime="00:05:14.61" resultid="1635" heatid="2404" lane="5" entrytime="00:05:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.60" />
                    <SPLIT distance="100" swimtime="00:01:08.01" />
                    <SPLIT distance="150" swimtime="00:01:47.54" />
                    <SPLIT distance="200" swimtime="00:02:26.64" />
                    <SPLIT distance="250" swimtime="00:03:12.85" />
                    <SPLIT distance="300" swimtime="00:04:01.24" />
                    <SPLIT distance="350" swimtime="00:04:38.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="438" swimtime="00:01:03.61" resultid="1636" heatid="2411" lane="6" entrytime="00:01:05.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carol" lastname="Nalle Bejes" birthdate="2010-04-20" gender="F" nation="BRA" license="377315" athleteid="1695" externalid="377315">
              <RESULTS>
                <RESULT eventid="1191" points="413" swimtime="00:00:38.07" resultid="1696" heatid="2380" lane="3" entrytime="00:00:38.25" entrycourse="SCM" />
                <RESULT eventid="1232" points="485" swimtime="00:02:51.24" resultid="1697" heatid="2386" lane="5" entrytime="00:03:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.21" />
                    <SPLIT distance="100" swimtime="00:01:22.84" />
                    <SPLIT distance="150" swimtime="00:02:06.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1444" points="440" swimtime="00:01:21.94" resultid="1698" heatid="2421" lane="8" entrytime="00:01:25.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" status="RJC" swimtime="00:00:00.00" resultid="1699" entrytime="00:02:55.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luana" lastname="Yoshie Kimura" birthdate="2010-07-08" gender="F" nation="BRA" license="391142" athleteid="1976" externalid="391142">
              <RESULTS>
                <RESULT eventid="1087" status="RJC" swimtime="00:00:00.00" resultid="1977" entrytime="00:02:53.29" entrycourse="SCM" />
                <RESULT eventid="1191" points="475" swimtime="00:00:36.35" resultid="1978" heatid="2380" lane="5" entrytime="00:00:37.92" entrycourse="SCM" />
                <RESULT eventid="1232" points="485" swimtime="00:02:51.18" resultid="1979" heatid="2386" lane="4" entrytime="00:03:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                    <SPLIT distance="100" swimtime="00:01:21.92" />
                    <SPLIT distance="150" swimtime="00:02:07.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="384" swimtime="00:05:56.11" resultid="1980" heatid="2403" lane="8" entrytime="00:06:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.28" />
                    <SPLIT distance="100" swimtime="00:01:24.58" />
                    <SPLIT distance="150" swimtime="00:02:12.19" />
                    <SPLIT distance="200" swimtime="00:02:59.17" />
                    <SPLIT distance="250" swimtime="00:03:43.69" />
                    <SPLIT distance="300" swimtime="00:04:30.89" />
                    <SPLIT distance="350" swimtime="00:05:14.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1444" points="499" swimtime="00:01:18.59" resultid="1981" heatid="2421" lane="3" entrytime="00:01:22.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Krupacz" birthdate="2008-04-18" gender="F" nation="BRA" license="329187" athleteid="1637" externalid="329187">
              <RESULTS>
                <RESULT eventid="1113" points="589" swimtime="00:00:30.12" resultid="1638" heatid="2367" lane="4" entrytime="00:00:30.70" entrycourse="SCM" />
                <RESULT eventid="1284" points="576" swimtime="00:02:22.94" resultid="1639" heatid="2396" lane="4" entrytime="00:02:25.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.84" />
                    <SPLIT distance="100" swimtime="00:01:08.36" />
                    <SPLIT distance="150" swimtime="00:01:45.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="583" swimtime="00:01:05.68" resultid="1640" heatid="2409" lane="4" entrytime="00:01:06.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Liz Skowronski" birthdate="2008-01-24" gender="F" nation="BRA" license="358245" athleteid="1718" externalid="358245">
              <RESULTS>
                <RESULT eventid="1113" points="346" swimtime="00:00:35.95" resultid="1719" heatid="2366" lane="4" entrytime="00:00:36.76" entrycourse="SCM" />
                <RESULT eventid="1284" points="377" swimtime="00:02:44.61" resultid="1720" heatid="2395" lane="4" entrytime="00:02:47.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.42" />
                    <SPLIT distance="100" swimtime="00:01:19.65" />
                    <SPLIT distance="150" swimtime="00:02:02.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="353" swimtime="00:01:17.62" resultid="1721" heatid="2408" lane="3" entrytime="00:01:17.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Blansky Hagebock" birthdate="2008-08-15" gender="M" nation="BRA" license="339123" athleteid="1688" externalid="339123">
              <RESULTS>
                <RESULT eventid="1126" points="530" swimtime="00:00:55.40" resultid="1689" heatid="2370" lane="7" entrytime="00:00:56.08" entrycourse="SCM" />
                <RESULT eventid="1405" points="451" swimtime="00:02:09.57" resultid="1690" heatid="2414" lane="6" entrytime="00:02:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                    <SPLIT distance="100" swimtime="00:01:02.78" />
                    <SPLIT distance="150" swimtime="00:01:36.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jennifer" lastname="De Abreu" birthdate="2009-11-07" gender="F" nation="BRA" license="356212" athleteid="1742" externalid="356212">
              <RESULTS>
                <RESULT eventid="1139" points="493" swimtime="00:01:03.60" resultid="1743" heatid="2372" lane="5" entrytime="00:01:03.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1061" points="459" swimtime="00:19:37.08" resultid="1744" heatid="2358" lane="5" entrytime="00:23:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                    <SPLIT distance="100" swimtime="00:01:13.06" />
                    <SPLIT distance="150" swimtime="00:01:52.32" />
                    <SPLIT distance="200" swimtime="00:02:30.69" />
                    <SPLIT distance="250" swimtime="00:03:09.65" />
                    <SPLIT distance="300" swimtime="00:03:49.26" />
                    <SPLIT distance="350" swimtime="00:04:28.20" />
                    <SPLIT distance="400" swimtime="00:05:07.15" />
                    <SPLIT distance="450" swimtime="00:05:46.20" />
                    <SPLIT distance="500" swimtime="00:06:25.60" />
                    <SPLIT distance="550" swimtime="00:07:05.24" />
                    <SPLIT distance="600" swimtime="00:07:44.22" />
                    <SPLIT distance="650" swimtime="00:08:22.34" />
                    <SPLIT distance="700" swimtime="00:09:02.13" />
                    <SPLIT distance="750" swimtime="00:09:42.27" />
                    <SPLIT distance="800" swimtime="00:10:21.73" />
                    <SPLIT distance="850" swimtime="00:11:01.49" />
                    <SPLIT distance="900" swimtime="00:11:41.82" />
                    <SPLIT distance="950" swimtime="00:12:22.13" />
                    <SPLIT distance="1000" swimtime="00:13:01.27" />
                    <SPLIT distance="1050" swimtime="00:13:40.59" />
                    <SPLIT distance="1100" swimtime="00:14:20.38" />
                    <SPLIT distance="1150" swimtime="00:15:01.06" />
                    <SPLIT distance="1200" swimtime="00:15:41.21" />
                    <SPLIT distance="1250" swimtime="00:16:21.20" />
                    <SPLIT distance="1300" swimtime="00:17:01.78" />
                    <SPLIT distance="1350" swimtime="00:17:41.11" />
                    <SPLIT distance="1400" swimtime="00:18:20.03" />
                    <SPLIT distance="1450" swimtime="00:18:57.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="395" swimtime="00:01:13.64" resultid="1745" heatid="2400" lane="6" entrytime="00:01:16.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="477" swimtime="00:02:21.10" resultid="1746" heatid="2412" lane="4" entrytime="00:02:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                    <SPLIT distance="100" swimtime="00:01:09.34" />
                    <SPLIT distance="150" swimtime="00:01:45.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolas" lastname="Mingorance Martins" birthdate="2007-10-13" gender="M" nation="BRA" license="393920" athleteid="1739" externalid="393920">
              <RESULTS>
                <RESULT eventid="1349" points="363" swimtime="00:05:28.96" resultid="1740" heatid="2404" lane="4" entrytime="00:05:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                    <SPLIT distance="100" swimtime="00:01:12.64" />
                    <SPLIT distance="150" swimtime="00:01:56.02" />
                    <SPLIT distance="200" swimtime="00:02:37.31" />
                    <SPLIT distance="250" swimtime="00:03:25.40" />
                    <SPLIT distance="300" swimtime="00:04:15.06" />
                    <SPLIT distance="350" swimtime="00:04:53.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="405" swimtime="00:09:55.14" resultid="1741" heatid="2425" lane="6" entrytime="00:12:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                    <SPLIT distance="100" swimtime="00:01:05.82" />
                    <SPLIT distance="150" swimtime="00:01:40.48" />
                    <SPLIT distance="200" swimtime="00:02:16.77" />
                    <SPLIT distance="250" swimtime="00:02:53.19" />
                    <SPLIT distance="300" swimtime="00:03:29.80" />
                    <SPLIT distance="350" swimtime="00:04:07.46" />
                    <SPLIT distance="400" swimtime="00:04:45.86" />
                    <SPLIT distance="450" swimtime="00:05:24.94" />
                    <SPLIT distance="500" swimtime="00:06:04.22" />
                    <SPLIT distance="550" swimtime="00:06:44.15" />
                    <SPLIT distance="600" swimtime="00:07:23.54" />
                    <SPLIT distance="650" swimtime="00:08:02.83" />
                    <SPLIT distance="700" swimtime="00:08:41.27" />
                    <SPLIT distance="750" swimtime="00:09:17.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Rodrigues Galvao" birthdate="2007-04-19" gender="M" nation="BRA" license="376586" athleteid="1677" externalid="376586">
              <RESULTS>
                <RESULT eventid="1271" points="471" swimtime="00:00:25.91" resultid="1678" heatid="2394" lane="6" entrytime="00:00:25.48" entrycourse="SCM" />
                <RESULT eventid="1431" points="514" swimtime="00:00:27.15" resultid="1679" heatid="2419" lane="4" entrytime="00:00:27.06" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Da Costa Riekes" birthdate="2008-06-19" gender="F" nation="BRA" license="331686" athleteid="1708" externalid="331686" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1139" points="513" swimtime="00:01:02.75" resultid="1709" heatid="2372" lane="3" entrytime="00:01:03.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="418" swimtime="00:01:12.26" resultid="1710" heatid="2400" lane="2" entrytime="00:01:16.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="514" swimtime="00:00:28.62" resultid="1711" heatid="2391" lane="5" entrytime="00:00:29.55" entrycourse="SCM" />
                <RESULT eventid="1418" points="473" swimtime="00:00:31.29" resultid="1712" heatid="2417" lane="4" entrytime="00:00:31.82" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="David Cella" birthdate="2008-02-17" gender="M" nation="BRA" license="341107" swrid="5634581" athleteid="1663" externalid="341107">
              <RESULTS>
                <RESULT eventid="1100" status="RJC" swimtime="00:00:00.00" resultid="1664" />
                <RESULT eventid="1271" points="589" swimtime="00:00:24.04" resultid="1665" heatid="2394" lane="4" entrytime="00:00:24.55" entrycourse="SCM" />
                <RESULT eventid="1126" points="612" swimtime="00:00:52.80" resultid="2350" heatid="2370" lane="6" entrytime="00:00:54.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="567" swimtime="00:00:30.13" resultid="2351" heatid="2378" lane="4" entrytime="00:00:30.47" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="De Krinski" birthdate="2007-07-20" gender="M" nation="BRA" license="334494" athleteid="1671" externalid="334494">
              <RESULTS>
                <RESULT eventid="1100" points="451" swimtime="00:00:28.82" resultid="1672" heatid="2365" lane="4" entrytime="00:00:28.27" entrycourse="SCM" />
                <RESULT eventid="1297" points="494" swimtime="00:02:13.58" resultid="1673" heatid="2398" lane="8" entrytime="00:02:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                    <SPLIT distance="100" swimtime="00:01:05.07" />
                    <SPLIT distance="150" swimtime="00:01:39.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" status="SICK" swimtime="00:00:00.00" resultid="1674" heatid="2411" lane="5" entrytime="00:01:00.21" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Bulla Lanaro" birthdate="2009-08-28" gender="F" nation="BRA" license="344301" athleteid="1651" externalid="344301">
              <RESULTS>
                <RESULT eventid="1139" points="550" swimtime="00:01:01.30" resultid="1652" heatid="2372" lane="4" entrytime="00:01:01.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="492" swimtime="00:02:31.50" resultid="1653" heatid="2376" lane="5" entrytime="00:02:29.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                    <SPLIT distance="100" swimtime="00:01:11.75" />
                    <SPLIT distance="150" swimtime="00:01:51.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="572" swimtime="00:01:05.09" resultid="1654" heatid="2400" lane="4" entrytime="00:01:05.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="552" swimtime="00:00:27.94" resultid="1655" heatid="2390" lane="4" entrytime="00:00:33.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabio" lastname="C Burak" birthdate="2009-08-29" gender="M" nation="BRA" license="343297" athleteid="1703" externalid="343297">
              <RESULTS>
                <RESULT eventid="1074" status="DSQ" swimtime="00:02:21.06" resultid="1704" heatid="2361" lane="1" entrytime="00:02:27.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                    <SPLIT distance="100" swimtime="00:01:08.37" />
                    <SPLIT distance="150" swimtime="00:01:47.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="426" swimtime="00:00:33.15" resultid="1705" heatid="2378" lane="2" entrytime="00:00:34.27" entrycourse="SCM" />
                <RESULT eventid="1245" points="397" swimtime="00:02:43.37" resultid="1706" heatid="2388" lane="3" entrytime="00:03:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.96" />
                    <SPLIT distance="100" swimtime="00:01:18.98" />
                    <SPLIT distance="150" swimtime="00:02:01.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="461" swimtime="00:01:11.51" resultid="1707" heatid="2424" lane="1" entrytime="00:01:12.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonia" lastname="Adam  Fracaro" birthdate="2010-04-27" gender="F" nation="BRA" license="382212" athleteid="1675" externalid="382212">
              <RESULTS>
                <RESULT eventid="1392" points="357" swimtime="00:02:35.39" resultid="1676" heatid="2412" lane="3" entrytime="00:02:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                    <SPLIT distance="100" swimtime="00:01:13.59" />
                    <SPLIT distance="150" swimtime="00:01:55.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Giuseppe Bulla Lanaro" birthdate="2007-05-22" gender="M" nation="BRA" license="331630" athleteid="1656" externalid="331630">
              <RESULTS>
                <RESULT eventid="1126" points="576" swimtime="00:00:53.88" resultid="1657" heatid="2370" lane="4" entrytime="00:00:53.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="593" swimtime="00:04:12.62" resultid="1658" heatid="2385" lane="5" entrytime="00:04:11.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.13" />
                    <SPLIT distance="100" swimtime="00:00:58.87" />
                    <SPLIT distance="150" swimtime="00:01:29.89" />
                    <SPLIT distance="200" swimtime="00:02:01.66" />
                    <SPLIT distance="250" swimtime="00:02:33.71" />
                    <SPLIT distance="300" swimtime="00:03:06.27" />
                    <SPLIT distance="350" swimtime="00:03:39.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="505" swimtime="00:00:25.30" resultid="1659" heatid="2394" lane="5" entrytime="00:00:24.91" entrycourse="SCM" />
                <RESULT eventid="1405" points="579" swimtime="00:01:59.16" resultid="1660" heatid="2415" lane="4" entrytime="00:01:56.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.16" />
                    <SPLIT distance="100" swimtime="00:00:56.84" />
                    <SPLIT distance="150" swimtime="00:01:28.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emily" lastname="Sayuri Tangueria De Lima" birthdate="2010-06-11" gender="F" nation="BRA" license="367215" athleteid="1691" externalid="367215">
              <RESULTS>
                <RESULT eventid="1165" points="358" swimtime="00:02:48.41" resultid="1692" heatid="2375" lane="3" entrytime="00:03:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                    <SPLIT distance="100" swimtime="00:01:17.39" />
                    <SPLIT distance="150" swimtime="00:02:02.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="466" swimtime="00:04:58.31" resultid="1693" heatid="2383" lane="1" entrytime="00:05:11.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.96" />
                    <SPLIT distance="100" swimtime="00:01:12.09" />
                    <SPLIT distance="150" swimtime="00:01:50.14" />
                    <SPLIT distance="200" swimtime="00:02:28.41" />
                    <SPLIT distance="250" swimtime="00:03:06.81" />
                    <SPLIT distance="300" swimtime="00:03:45.37" />
                    <SPLIT distance="350" swimtime="00:04:22.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1418" points="364" swimtime="00:00:34.13" resultid="1694" heatid="2417" lane="1" entrytime="00:00:34.01" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Garcia De Fraga" birthdate="2009-03-24" gender="M" nation="BRA" license="342147" athleteid="1641" externalid="342147" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1074" points="504" swimtime="00:02:17.69" resultid="1642" heatid="2361" lane="4" entrytime="00:02:11.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                    <SPLIT distance="100" swimtime="00:01:04.23" />
                    <SPLIT distance="150" swimtime="00:01:44.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="442" swimtime="00:00:29.01" resultid="1643" heatid="2365" lane="8" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1323" points="480" swimtime="00:01:01.01" resultid="1644" heatid="2401" lane="2" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="491" swimtime="00:01:01.26" resultid="1645" heatid="2411" lane="4" entrytime="00:00:59.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benito" lastname="Alves Sant&apos;Ana" birthdate="2009-06-01" gender="M" nation="BRA" license="376585" athleteid="1722" externalid="376585">
              <RESULTS>
                <RESULT eventid="1219" points="525" swimtime="00:04:22.96" resultid="1723" heatid="2385" lane="2" entrytime="00:04:27.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.67" />
                    <SPLIT distance="100" swimtime="00:01:01.67" />
                    <SPLIT distance="150" swimtime="00:01:34.23" />
                    <SPLIT distance="200" swimtime="00:02:07.51" />
                    <SPLIT distance="250" swimtime="00:02:41.62" />
                    <SPLIT distance="300" swimtime="00:03:15.54" />
                    <SPLIT distance="350" swimtime="00:03:50.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="478" swimtime="00:05:00.22" resultid="1724" heatid="2404" lane="3" entrytime="00:05:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.16" />
                    <SPLIT distance="100" swimtime="00:01:09.36" />
                    <SPLIT distance="150" swimtime="00:01:46.47" />
                    <SPLIT distance="200" swimtime="00:02:23.88" />
                    <SPLIT distance="250" swimtime="00:03:07.92" />
                    <SPLIT distance="300" swimtime="00:03:52.07" />
                    <SPLIT distance="350" swimtime="00:04:27.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="541" swimtime="00:09:00.29" resultid="1725" heatid="2426" lane="2" entrytime="00:09:05.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                    <SPLIT distance="100" swimtime="00:01:04.11" />
                    <SPLIT distance="150" swimtime="00:01:38.54" />
                    <SPLIT distance="200" swimtime="00:02:11.78" />
                    <SPLIT distance="250" swimtime="00:02:45.89" />
                    <SPLIT distance="300" swimtime="00:03:19.73" />
                    <SPLIT distance="350" swimtime="00:03:53.88" />
                    <SPLIT distance="400" swimtime="00:04:28.65" />
                    <SPLIT distance="450" swimtime="00:05:03.29" />
                    <SPLIT distance="500" swimtime="00:05:37.55" />
                    <SPLIT distance="550" swimtime="00:06:11.90" />
                    <SPLIT distance="600" swimtime="00:06:45.64" />
                    <SPLIT distance="650" swimtime="00:07:20.42" />
                    <SPLIT distance="700" swimtime="00:07:54.83" />
                    <SPLIT distance="750" swimtime="00:08:28.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Braga" birthdate="2010-05-07" gender="M" nation="BRA" license="378345" athleteid="1629" externalid="378345">
              <RESULTS>
                <RESULT eventid="1245" points="429" swimtime="00:02:39.26" resultid="1630" heatid="2389" lane="6" entrytime="00:02:40.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                    <SPLIT distance="100" swimtime="00:01:14.67" />
                    <SPLIT distance="150" swimtime="00:01:56.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="426" swimtime="00:01:13.45" resultid="1631" heatid="2424" lane="7" entrytime="00:01:12.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Daniele Silva" birthdate="2010-07-06" gender="F" nation="BRA" license="359593" athleteid="1730" externalid="359593" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1113" points="408" swimtime="00:00:34.03" resultid="1731" heatid="2367" lane="7" entrytime="00:00:34.61" entrycourse="SCM" />
                <RESULT eventid="1284" points="416" swimtime="00:02:39.22" resultid="1732" heatid="2395" lane="2" entrytime="00:03:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.95" />
                    <SPLIT distance="100" swimtime="00:01:18.43" />
                    <SPLIT distance="150" swimtime="00:01:59.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="378" swimtime="00:01:15.90" resultid="1733" heatid="2409" lane="1" entrytime="00:01:15.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabrizio" lastname="Bulla Lanaro" birthdate="2009-08-28" gender="M" nation="BRA" license="344303" athleteid="1680" externalid="344303">
              <RESULTS>
                <RESULT eventid="1152" points="387" swimtime="00:02:26.52" resultid="1681" heatid="2373" lane="6" entrytime="00:03:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.78" />
                    <SPLIT distance="100" swimtime="00:01:08.53" />
                    <SPLIT distance="150" swimtime="00:01:47.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1323" points="446" swimtime="00:01:02.50" resultid="1682" heatid="2402" lane="1" entrytime="00:01:03.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="488" swimtime="00:00:27.61" resultid="1683" heatid="2419" lane="6" entrytime="00:00:28.28" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcus" lastname="Vinicius De Almeida" birthdate="2009-06-16" gender="M" nation="BRA" license="348099" athleteid="1726" externalid="348099">
              <RESULTS>
                <RESULT eventid="1178" points="448" swimtime="00:00:32.60" resultid="1727" heatid="2378" lane="3" entrytime="00:00:32.37" entrycourse="SCM" />
                <RESULT eventid="1245" points="473" swimtime="00:02:34.20" resultid="1728" heatid="2389" lane="3" entrytime="00:02:38.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                    <SPLIT distance="100" swimtime="00:01:13.21" />
                    <SPLIT distance="150" swimtime="00:01:54.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="525" swimtime="00:01:08.51" resultid="1729" heatid="2424" lane="3" entrytime="00:01:10.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Sieck" birthdate="2011-01-20" gender="F" nation="BRA" license="382234" athleteid="1734" externalid="382234">
              <RESULTS>
                <RESULT comment=" (Horário: 10:00)" eventid="1418" status="DSQ" swimtime="00:00:42.26" resultid="1735" heatid="2416" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Inoue Kuroda" birthdate="2009-04-18" gender="M" nation="BRA" license="324700" athleteid="1684" externalid="324700">
              <RESULTS>
                <RESULT eventid="1297" points="405" swimtime="00:02:22.75" resultid="1685" heatid="2397" lane="3" entrytime="00:02:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.91" />
                    <SPLIT distance="100" swimtime="00:01:07.23" />
                    <SPLIT distance="150" swimtime="00:01:44.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="447" swimtime="00:09:36.03" resultid="1686" heatid="2426" lane="6" entrytime="00:09:03.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.85" />
                    <SPLIT distance="100" swimtime="00:01:05.90" />
                    <SPLIT distance="150" swimtime="00:01:40.65" />
                    <SPLIT distance="200" swimtime="00:02:15.47" />
                    <SPLIT distance="250" swimtime="00:02:50.46" />
                    <SPLIT distance="300" swimtime="00:03:27.29" />
                    <SPLIT distance="350" swimtime="00:04:04.55" />
                    <SPLIT distance="400" swimtime="00:04:41.96" />
                    <SPLIT distance="450" swimtime="00:05:19.67" />
                    <SPLIT distance="500" swimtime="00:05:57.76" />
                    <SPLIT distance="550" swimtime="00:06:35.63" />
                    <SPLIT distance="600" swimtime="00:07:13.06" />
                    <SPLIT distance="650" swimtime="00:07:51.64" />
                    <SPLIT distance="700" swimtime="00:08:29.15" />
                    <SPLIT distance="750" swimtime="00:09:06.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1405" points="512" swimtime="00:02:04.17" resultid="1687" heatid="2414" lane="1" entrytime="00:02:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.16" />
                    <SPLIT distance="100" swimtime="00:00:59.86" />
                    <SPLIT distance="150" swimtime="00:01:32.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Fernandes" birthdate="2010-03-13" gender="M" nation="BRA" license="339266" athleteid="1661" externalid="339266">
              <RESULTS>
                <RESULT eventid="1297" points="392" swimtime="00:02:24.24" resultid="1662" heatid="2397" lane="4" entrytime="00:02:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.06" />
                    <SPLIT distance="100" swimtime="00:01:09.90" />
                    <SPLIT distance="150" swimtime="00:01:46.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1364" points="603" swimtime="00:03:36.27" resultid="1749" heatid="2407" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.99" />
                    <SPLIT distance="100" swimtime="00:00:53.10" />
                    <SPLIT distance="150" swimtime="00:01:18.98" />
                    <SPLIT distance="200" swimtime="00:01:47.63" />
                    <SPLIT distance="250" swimtime="00:02:14.18" />
                    <SPLIT distance="300" swimtime="00:02:43.18" />
                    <SPLIT distance="350" swimtime="00:03:08.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1663" number="1" />
                    <RELAYPOSITION athleteid="1688" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1677" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1656" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1485" status="DSQ" swimtime="00:04:04.16" resultid="1750" heatid="2428" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.80" />
                    <SPLIT distance="100" swimtime="00:01:01.13" />
                    <SPLIT distance="150" swimtime="00:01:33.26" />
                    <SPLIT distance="200" swimtime="00:02:09.58" />
                    <SPLIT distance="250" swimtime="00:02:37.57" />
                    <SPLIT distance="300" swimtime="00:03:11.25" />
                    <SPLIT distance="350" swimtime="00:03:35.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1641" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="1726" number="2" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION athleteid="1680" number="3" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION athleteid="1663" number="4" reactiontime="0" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1362" points="557" swimtime="00:04:09.67" resultid="1747" heatid="2406" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.39" />
                    <SPLIT distance="100" swimtime="00:01:01.05" />
                    <SPLIT distance="150" swimtime="00:01:30.87" />
                    <SPLIT distance="200" swimtime="00:02:05.00" />
                    <SPLIT distance="250" swimtime="00:02:34.75" />
                    <SPLIT distance="300" swimtime="00:03:07.69" />
                    <SPLIT distance="350" swimtime="00:03:37.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1651" number="1" />
                    <RELAYPOSITION athleteid="1730" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1742" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1708" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1483" points="544" swimtime="00:04:34.82" resultid="1748" heatid="2427" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                    <SPLIT distance="100" swimtime="00:01:05.95" />
                    <SPLIT distance="150" swimtime="00:01:43.34" />
                    <SPLIT distance="200" swimtime="00:02:25.27" />
                    <SPLIT distance="250" swimtime="00:02:56.67" />
                    <SPLIT distance="300" swimtime="00:03:32.64" />
                    <SPLIT distance="350" swimtime="00:04:02.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1637" number="1" />
                    <RELAYPOSITION athleteid="1976" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1651" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1708" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1204" status="DSQ" swimtime="00:01:55.58" resultid="1751" heatid="2381" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                    <SPLIT distance="100" swimtime="00:01:00.93" />
                    <SPLIT distance="150" swimtime="00:01:30.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1637" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="1663" number="2" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION athleteid="1651" number="3" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION athleteid="1656" number="4" reactiontime="0" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="1490" nation="BRA" region="PR" clubid="1982" name="Seleção De Ponta Grossa/PR" shortname="Ponta Grossa">
          <ATHLETES>
            <ATHLETE firstname="Gabriela" lastname="Lievore" birthdate="2010-06-07" gender="F" nation="BRA" license="414856" athleteid="2033" externalid="414856">
              <RESULTS>
                <RESULT eventid="1139" points="290" swimtime="00:01:15.89" resultid="2034" heatid="2371" lane="2" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" status="DNS" swimtime="00:00:00.00" resultid="2035" heatid="2379" lane="1" />
                <RESULT eventid="1258" points="317" swimtime="00:00:33.62" resultid="2036" heatid="2390" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Brenda" lastname="Gabriele Carvalho" birthdate="2010-04-11" gender="F" nation="BRA" license="399557" athleteid="2021" externalid="399557">
              <RESULTS>
                <RESULT eventid="1087" points="256" swimtime="00:03:11.77" resultid="2022" heatid="2362" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.89" />
                    <SPLIT distance="150" swimtime="00:02:28.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="244" swimtime="00:01:27.78" resultid="2023" heatid="2408" lane="1" entrytime="00:01:31.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Reda" birthdate="2007-05-21" gender="F" nation="BRA" license="316228" athleteid="1998" externalid="316228">
              <RESULTS>
                <RESULT eventid="1139" status="WDR" swimtime="00:00:00.00" resultid="1999" entrytime="00:01:15.00" entrycourse="SCM" />
                <RESULT eventid="1113" status="WDR" swimtime="00:00:00.00" resultid="2000" entrytime="00:00:40.00" entrycourse="SCM" />
                <RESULT eventid="1258" status="WDR" swimtime="00:00:00.00" resultid="2001" entrytime="00:00:33.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Chi Kravchychyn" birthdate="2009-09-27" gender="M" nation="BRA" license="344268" athleteid="1988" externalid="344268">
              <RESULTS>
                <RESULT eventid="1152" points="371" swimtime="00:02:28.58" resultid="1989" heatid="2373" lane="4" entrytime="00:03:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.86" />
                    <SPLIT distance="100" swimtime="00:01:07.64" />
                    <SPLIT distance="150" swimtime="00:01:46.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1245" points="521" swimtime="00:02:29.29" resultid="1990" heatid="2389" lane="5" entrytime="00:02:29.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                    <SPLIT distance="100" swimtime="00:01:12.95" />
                    <SPLIT distance="150" swimtime="00:01:51.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="455" swimtime="00:05:05.17" resultid="1991" heatid="2405" lane="6" entrytime="00:04:59.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                    <SPLIT distance="100" swimtime="00:01:09.20" />
                    <SPLIT distance="150" swimtime="00:01:50.54" />
                    <SPLIT distance="200" swimtime="00:02:30.63" />
                    <SPLIT distance="250" swimtime="00:03:13.42" />
                    <SPLIT distance="300" swimtime="00:03:56.81" />
                    <SPLIT distance="350" swimtime="00:04:31.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="480" swimtime="00:01:10.60" resultid="1992" heatid="2424" lane="5" entrytime="00:01:09.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Carraro Borges" birthdate="2009-05-11" gender="M" nation="BRA" license="345590" athleteid="2016" externalid="345590" level="SAGRADA FA">
              <RESULTS>
                <RESULT eventid="1126" points="412" swimtime="00:01:00.25" resultid="2017" heatid="2368" lane="4" entrytime="00:01:06.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="425" swimtime="00:04:42.20" resultid="2018" heatid="2384" lane="4" entrytime="00:04:44.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.53" />
                    <SPLIT distance="100" swimtime="00:01:06.91" />
                    <SPLIT distance="150" swimtime="00:01:42.62" />
                    <SPLIT distance="200" swimtime="00:02:19.16" />
                    <SPLIT distance="250" swimtime="00:02:55.39" />
                    <SPLIT distance="300" swimtime="00:03:32.02" />
                    <SPLIT distance="350" swimtime="00:04:07.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="371" swimtime="00:10:12.86" resultid="2019" heatid="2426" lane="8" entrytime="00:10:05.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="100" swimtime="00:01:11.43" />
                    <SPLIT distance="150" swimtime="00:01:49.93" />
                    <SPLIT distance="200" swimtime="00:02:28.46" />
                    <SPLIT distance="250" swimtime="00:03:07.48" />
                    <SPLIT distance="300" swimtime="00:03:46.54" />
                    <SPLIT distance="350" swimtime="00:04:25.49" />
                    <SPLIT distance="400" swimtime="00:05:04.82" />
                    <SPLIT distance="450" swimtime="00:05:44.56" />
                    <SPLIT distance="500" swimtime="00:06:22.60" />
                    <SPLIT distance="550" swimtime="00:07:01.19" />
                    <SPLIT distance="600" swimtime="00:07:39.19" />
                    <SPLIT distance="650" swimtime="00:08:18.08" />
                    <SPLIT distance="700" swimtime="00:08:56.49" />
                    <SPLIT distance="750" swimtime="00:09:34.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1405" points="406" swimtime="00:02:14.16" resultid="2020" heatid="2414" lane="2" entrytime="00:02:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.36" />
                    <SPLIT distance="100" swimtime="00:01:05.15" />
                    <SPLIT distance="150" swimtime="00:01:39.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Barbara" lastname="Campagnoli" birthdate="2009-04-13" gender="F" nation="BRA" license="366915" athleteid="1993" externalid="366915">
              <RESULTS>
                <RESULT eventid="1139" points="509" swimtime="00:01:02.92" resultid="1994" heatid="2372" lane="6" entrytime="00:01:04.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="501" swimtime="00:00:31.78" resultid="1995" heatid="2367" lane="5" entrytime="00:00:32.73" entrycourse="SCM" />
                <RESULT eventid="1284" points="432" swimtime="00:02:37.22" resultid="1996" heatid="2395" lane="6" entrytime="00:03:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                    <SPLIT distance="100" swimtime="00:01:15.63" />
                    <SPLIT distance="150" swimtime="00:01:57.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="418" swimtime="00:01:13.36" resultid="1997" heatid="2409" lane="3" entrytime="00:01:13.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Gueiber Montes" birthdate="2009-03-09" gender="M" nation="BRA" license="342154" athleteid="1983" externalid="342154">
              <RESULTS>
                <RESULT eventid="1126" points="576" swimtime="00:00:53.88" resultid="1984" heatid="2370" lane="3" entrytime="00:00:54.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="562" swimtime="00:04:17.17" resultid="1985" heatid="2385" lane="7" entrytime="00:04:27.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                    <SPLIT distance="100" swimtime="00:01:02.30" />
                    <SPLIT distance="150" swimtime="00:01:36.05" />
                    <SPLIT distance="200" swimtime="00:02:09.12" />
                    <SPLIT distance="250" swimtime="00:02:42.52" />
                    <SPLIT distance="300" swimtime="00:03:15.58" />
                    <SPLIT distance="350" swimtime="00:03:46.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="493" swimtime="00:00:25.51" resultid="1986" heatid="2394" lane="3" entrytime="00:00:25.27" entrycourse="SCM" />
                <RESULT eventid="1405" points="581" swimtime="00:01:59.05" resultid="1987" heatid="2414" lane="5" entrytime="00:02:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.80" />
                    <SPLIT distance="100" swimtime="00:00:58.65" />
                    <SPLIT distance="150" swimtime="00:01:29.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Carolina Babiuki" birthdate="2007-02-06" gender="F" nation="BRA" license="316227" athleteid="2002" externalid="316227" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1113" status="WDR" swimtime="00:00:00.00" resultid="2003" entrytime="00:00:31.79" entrycourse="SCM" />
                <RESULT eventid="1284" status="WDR" swimtime="00:00:00.00" resultid="2004" entrytime="00:03:18.00" entrycourse="SCM" />
                <RESULT eventid="1258" status="WDR" swimtime="00:00:00.00" resultid="2005" entrytime="00:00:28.53" entrycourse="SCM" />
                <RESULT eventid="1366" status="WDR" swimtime="00:00:00.00" resultid="2006" entrytime="00:01:12.31" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Franca Berger" birthdate="2010-05-07" gender="F" nation="BRA" license="399692" athleteid="2029" externalid="399692">
              <RESULTS>
                <RESULT eventid="1191" points="279" swimtime="00:00:43.40" resultid="2030" heatid="2379" lane="3" entrytime="00:00:44.95" entrycourse="SCM" />
                <RESULT eventid="1444" points="232" swimtime="00:01:41.44" resultid="2031" heatid="2420" lane="2" entrytime="00:01:42.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1418" status="DNS" swimtime="00:00:00.00" resultid="2032" heatid="2416" lane="3" entrytime="00:00:47.55" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Delinski" birthdate="2009-11-28" gender="F" nation="BRA" license="385190" athleteid="2007" externalid="385190">
              <RESULTS>
                <RESULT eventid="1191" points="393" swimtime="00:00:38.70" resultid="2008" heatid="2379" lane="5" entrytime="00:00:41.86" entrycourse="SCM" />
                <RESULT eventid="1232" points="332" swimtime="00:03:14.25" resultid="2009" heatid="2387" lane="8" entrytime="00:03:32.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.13" />
                    <SPLIT distance="100" swimtime="00:01:34.09" />
                    <SPLIT distance="150" swimtime="00:02:24.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1444" points="406" swimtime="00:01:24.18" resultid="2010" heatid="2420" lane="3" entrytime="00:01:31.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Fegert" birthdate="2009-04-13" gender="M" nation="BRA" license="353813" athleteid="2011" externalid="353813">
              <RESULTS>
                <RESULT eventid="1126" points="468" swimtime="00:00:57.75" resultid="2012" heatid="2369" lane="8" entrytime="00:01:06.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1323" points="456" swimtime="00:01:02.05" resultid="2013" heatid="2401" lane="4" entrytime="00:01:05.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="457" swimtime="00:00:26.17" resultid="2014" heatid="2393" lane="5" entrytime="00:00:27.72" entrycourse="SCM" />
                <RESULT eventid="1431" points="444" swimtime="00:00:28.50" resultid="2015" heatid="2419" lane="2" entrytime="00:00:28.38" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Augusto" lastname="Tramontin" birthdate="2011-11-29" gender="M" nation="BRA" license="399691" athleteid="2024" externalid="399691">
              <RESULTS>
                <RESULT eventid="1100" points="269" swimtime="00:00:34.25" resultid="2025" heatid="2365" lane="1" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1178" points="363" swimtime="00:00:34.97" resultid="2026" heatid="2377" lane="3" entrytime="00:00:38.39" entrycourse="SCM" />
                <RESULT eventid="1271" points="345" swimtime="00:00:28.73" resultid="2027" heatid="2393" lane="1" entrytime="00:00:28.93" entrycourse="SCM" />
                <RESULT eventid="1457" points="340" swimtime="00:01:19.19" resultid="2028" heatid="2423" lane="7" entrytime="00:01:26.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="PONTA GROSSA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1364" points="490" swimtime="00:03:51.69" resultid="2039" heatid="2407" lane="3" entrytime="00:03:41.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.48" />
                    <SPLIT distance="100" swimtime="00:00:54.81" />
                    <SPLIT distance="150" swimtime="00:01:22.08" />
                    <SPLIT distance="200" swimtime="00:01:52.96" />
                    <SPLIT distance="250" swimtime="00:02:20.16" />
                    <SPLIT distance="300" swimtime="00:02:51.11" />
                    <SPLIT distance="350" swimtime="00:03:19.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1983" number="1" />
                    <RELAYPOSITION athleteid="1988" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2011" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="2016" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1485" status="DSQ" swimtime="00:04:16.21" resultid="2040" heatid="2428" lane="3" entrytime="00:04:09.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.43" />
                    <SPLIT distance="100" swimtime="00:01:01.41" />
                    <SPLIT distance="150" swimtime="00:01:34.38" />
                    <SPLIT distance="200" swimtime="00:02:12.51" />
                    <SPLIT distance="250" swimtime="00:02:41.21" />
                    <SPLIT distance="300" swimtime="00:03:15.03" />
                    <SPLIT distance="350" swimtime="00:03:43.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1983" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="1988" number="2" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION athleteid="2011" number="3" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION athleteid="2016" number="4" reactiontime="0" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="PONTA GROSSA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1362" points="325" swimtime="00:04:58.60" resultid="2037" heatid="2406" lane="5" entrytime="00:04:15.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                    <SPLIT distance="100" swimtime="00:01:05.29" />
                    <SPLIT distance="150" swimtime="00:01:42.17" />
                    <SPLIT distance="200" swimtime="00:02:24.98" />
                    <SPLIT distance="250" swimtime="00:03:00.19" />
                    <SPLIT distance="300" swimtime="00:03:41.93" />
                    <SPLIT distance="350" swimtime="00:04:17.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1993" number="1" />
                    <RELAYPOSITION athleteid="2021" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2033" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="2029" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1483" points="292" swimtime="00:05:37.87" resultid="2038" heatid="2427" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                    <SPLIT distance="100" swimtime="00:01:14.90" />
                    <SPLIT distance="150" swimtime="00:02:03.58" />
                    <SPLIT distance="200" swimtime="00:02:58.22" />
                    <SPLIT distance="250" swimtime="00:03:35.52" />
                    <SPLIT distance="300" swimtime="00:04:23.61" />
                    <SPLIT distance="350" swimtime="00:04:58.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1993" number="1" />
                    <RELAYPOSITION athleteid="2021" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2007" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="2033" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="PONTA GROSSA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1204" status="DSQ" swimtime="00:02:03.46" resultid="2041" heatid="2381" lane="6">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1993" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="2007" number="2" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION athleteid="1988" number="3" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION athleteid="1983" number="4" reactiontime="0" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="1488" nation="BRA" region="PR" clubid="1858" name="Seleção De Maringá/PR" shortname="Maringá">
          <ATHLETES>
            <ATHLETE firstname="Tiago" lastname="Ficher Delmont Pais" birthdate="2010-07-15" gender="M" nation="BRA" license="338533" athleteid="1869" externalid="338533">
              <RESULTS>
                <RESULT eventid="1152" points="335" swimtime="00:02:33.80" resultid="1870" heatid="2373" lane="3" entrytime="00:03:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                    <SPLIT distance="100" swimtime="00:01:12.92" />
                    <SPLIT distance="150" swimtime="00:01:54.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="378" swimtime="00:02:31.49" resultid="1871" heatid="2361" lane="2" entrytime="00:02:23.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.67" />
                    <SPLIT distance="100" swimtime="00:01:07.88" />
                    <SPLIT distance="150" swimtime="00:01:55.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1323" points="492" swimtime="00:01:00.52" resultid="1872" heatid="2402" lane="5" entrytime="00:01:01.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="518" swimtime="00:00:27.08" resultid="1873" heatid="2419" lane="5" entrytime="00:00:27.33" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Mochiutti Carneiro" birthdate="2010-04-22" gender="F" nation="BRA" license="370670" athleteid="1944" externalid="370670">
              <RESULTS>
                <RESULT eventid="1165" points="291" swimtime="00:03:00.47" resultid="1945" heatid="2376" lane="2" entrytime="00:02:54.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                    <SPLIT distance="100" swimtime="00:01:22.32" />
                    <SPLIT distance="150" swimtime="00:02:10.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="414" swimtime="00:05:10.26" resultid="1946" heatid="2383" lane="7" entrytime="00:05:08.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                    <SPLIT distance="100" swimtime="00:01:13.15" />
                    <SPLIT distance="150" swimtime="00:01:51.91" />
                    <SPLIT distance="200" swimtime="00:02:31.46" />
                    <SPLIT distance="250" swimtime="00:03:11.89" />
                    <SPLIT distance="300" swimtime="00:03:52.44" />
                    <SPLIT distance="350" swimtime="00:04:32.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="333" swimtime="00:06:13.46" resultid="1947" heatid="2403" lane="7" entrytime="00:06:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.29" />
                    <SPLIT distance="100" swimtime="00:01:25.25" />
                    <SPLIT distance="150" swimtime="00:02:16.04" />
                    <SPLIT distance="200" swimtime="00:03:05.09" />
                    <SPLIT distance="250" swimtime="00:03:59.27" />
                    <SPLIT distance="300" swimtime="00:04:53.80" />
                    <SPLIT distance="350" swimtime="00:05:34.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1418" points="388" swimtime="00:00:33.40" resultid="1948" heatid="2417" lane="5" entrytime="00:00:31.98" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wellington" lastname="De Lima" birthdate="2008-03-01" gender="M" nation="BRA" license="370024" athleteid="1874" externalid="370024">
              <RESULTS>
                <RESULT eventid="1126" points="446" swimtime="00:00:58.66" resultid="1875" heatid="2370" lane="1" entrytime="00:00:56.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="390" swimtime="00:00:30.25" resultid="1876" heatid="2365" lane="5" entrytime="00:00:30.29" entrycourse="SCM" />
                <RESULT eventid="1271" points="473" swimtime="00:00:25.87" resultid="1877" heatid="2394" lane="7" entrytime="00:00:25.99" entrycourse="SCM" />
                <RESULT eventid="1379" points="363" swimtime="00:01:07.74" resultid="1878" heatid="2411" lane="7" entrytime="00:01:06.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Henrique Goes" birthdate="2008-10-26" gender="M" nation="BRA" license="392105" athleteid="1960" externalid="392105">
              <RESULTS>
                <RESULT eventid="1470" points="268" swimtime="00:11:22.92" resultid="1961" heatid="2425" lane="3" entrytime="00:11:32.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.10" />
                    <SPLIT distance="100" swimtime="00:01:16.72" />
                    <SPLIT distance="150" swimtime="00:01:59.38" />
                    <SPLIT distance="200" swimtime="00:02:42.85" />
                    <SPLIT distance="250" swimtime="00:03:26.49" />
                    <SPLIT distance="300" swimtime="00:04:10.09" />
                    <SPLIT distance="350" swimtime="00:04:54.33" />
                    <SPLIT distance="400" swimtime="00:05:38.49" />
                    <SPLIT distance="450" swimtime="00:06:22.51" />
                    <SPLIT distance="500" swimtime="00:07:06.57" />
                    <SPLIT distance="550" swimtime="00:07:50.39" />
                    <SPLIT distance="600" swimtime="00:08:33.82" />
                    <SPLIT distance="650" swimtime="00:09:16.85" />
                    <SPLIT distance="700" swimtime="00:09:59.85" />
                    <SPLIT distance="750" swimtime="00:10:42.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Batista Sanchez" birthdate="2009-05-22" gender="M" nation="BRA" license="370668" athleteid="1879" externalid="370668">
              <RESULTS>
                <RESULT eventid="1178" points="365" swimtime="00:00:34.89" resultid="1880" heatid="2378" lane="7" entrytime="00:00:34.30" entrycourse="SCM" />
                <RESULT eventid="1245" points="395" swimtime="00:02:43.67" resultid="1881" heatid="2389" lane="7" entrytime="00:02:41.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.68" />
                    <SPLIT distance="100" swimtime="00:01:17.89" />
                    <SPLIT distance="150" swimtime="00:02:00.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="350" swimtime="00:05:33.07" resultid="1882" heatid="2405" lane="8" entrytime="00:05:48.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.35" />
                    <SPLIT distance="100" swimtime="00:01:14.48" />
                    <SPLIT distance="150" swimtime="00:02:00.92" />
                    <SPLIT distance="200" swimtime="00:02:46.58" />
                    <SPLIT distance="250" swimtime="00:03:30.91" />
                    <SPLIT distance="300" swimtime="00:04:16.31" />
                    <SPLIT distance="350" swimtime="00:04:55.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="410" swimtime="00:01:14.41" resultid="1883" heatid="2424" lane="2" entrytime="00:01:11.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Otavio Costa" birthdate="2009-01-28" gender="M" nation="BRA" license="370666" athleteid="1937" externalid="370666">
              <RESULTS>
                <RESULT eventid="1074" points="280" swimtime="00:02:47.53" resultid="1938" heatid="2360" lane="6" entrytime="00:02:49.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                    <SPLIT distance="100" swimtime="00:01:24.04" />
                    <SPLIT distance="150" swimtime="00:02:10.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carina" lastname="Costa Profeta" birthdate="2008-03-20" gender="F" nation="BRA" license="366964" athleteid="1895" externalid="366964">
              <RESULTS>
                <RESULT eventid="1087" points="412" swimtime="00:02:43.68" resultid="1896" heatid="2363" lane="3" entrytime="00:02:41.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.22" />
                    <SPLIT distance="100" swimtime="00:01:16.68" />
                    <SPLIT distance="150" swimtime="00:02:01.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="464" swimtime="00:00:36.62" resultid="1897" heatid="2380" lane="4" entrytime="00:00:35.68" entrycourse="SCM" />
                <RESULT eventid="1232" points="457" swimtime="00:02:54.64" resultid="1898" heatid="2387" lane="3" entrytime="00:03:00.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.80" />
                    <SPLIT distance="100" swimtime="00:01:22.75" />
                    <SPLIT distance="150" swimtime="00:02:08.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1444" points="486" swimtime="00:01:19.31" resultid="1899" heatid="2421" lane="5" entrytime="00:01:20.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Casavechia Carraro" birthdate="2009-07-28" gender="M" nation="BRA" license="368150" athleteid="1864" externalid="368150">
              <RESULTS>
                <RESULT eventid="1126" points="629" swimtime="00:00:52.32" resultid="1865" heatid="2370" lane="5" entrytime="00:00:54.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1323" points="535" swimtime="00:00:58.82" resultid="1866" heatid="2402" lane="4" entrytime="00:00:59.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="536" swimtime="00:04:21.17" resultid="1867" heatid="2385" lane="6" entrytime="00:04:24.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.00" />
                    <SPLIT distance="100" swimtime="00:01:01.64" />
                    <SPLIT distance="150" swimtime="00:01:35.48" />
                    <SPLIT distance="200" swimtime="00:02:09.20" />
                    <SPLIT distance="250" swimtime="00:02:42.77" />
                    <SPLIT distance="300" swimtime="00:03:16.12" />
                    <SPLIT distance="350" swimtime="00:03:48.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1405" status="DSQ" swimtime="00:01:57.32" resultid="1868" heatid="2415" lane="5" entrytime="00:02:00.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                    <SPLIT distance="100" swimtime="00:00:56.93" />
                    <SPLIT distance="150" swimtime="00:01:27.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Antonio Mendes" birthdate="2008-12-04" gender="M" nation="BRA" license="366962" athleteid="1910" externalid="366962">
              <RESULTS>
                <RESULT eventid="1074" points="445" swimtime="00:02:23.51" resultid="1911" heatid="2361" lane="7" entrytime="00:02:25.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.86" />
                    <SPLIT distance="100" swimtime="00:01:08.41" />
                    <SPLIT distance="150" swimtime="00:01:47.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="505" swimtime="00:00:31.32" resultid="1912" heatid="2378" lane="5" entrytime="00:00:31.32" entrycourse="SCM" />
                <RESULT eventid="1245" points="512" swimtime="00:02:30.17" resultid="1913" heatid="2389" lane="4" entrytime="00:02:28.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                    <SPLIT distance="100" swimtime="00:01:11.97" />
                    <SPLIT distance="150" swimtime="00:01:51.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="503" swimtime="00:01:09.50" resultid="1914" heatid="2424" lane="4" entrytime="00:01:08.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Ghelere" birthdate="2011-04-03" gender="F" nation="BRA" license="368146" athleteid="1930" externalid="368146">
              <RESULTS>
                <RESULT eventid="1087" points="245" swimtime="00:03:14.67" resultid="1931" heatid="2363" lane="1" entrytime="00:03:12.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                    <SPLIT distance="100" swimtime="00:01:26.91" />
                    <SPLIT distance="150" swimtime="00:02:30.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="305" swimtime="00:02:43.75" resultid="1932" heatid="2413" lane="8" entrytime="00:02:41.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                    <SPLIT distance="100" swimtime="00:01:19.13" />
                    <SPLIT distance="150" swimtime="00:02:02.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Garcia Cavalcante" birthdate="2008-08-11" gender="M" nation="BRA" license="369676" swrid="5603841" athleteid="1884" externalid="369676">
              <RESULTS>
                <RESULT eventid="1219" points="407" swimtime="00:04:46.27" resultid="1885" heatid="2385" lane="8" entrytime="00:04:43.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                    <SPLIT distance="100" swimtime="00:01:06.99" />
                    <SPLIT distance="150" swimtime="00:01:43.73" />
                    <SPLIT distance="200" swimtime="00:02:20.25" />
                    <SPLIT distance="250" swimtime="00:02:56.30" />
                    <SPLIT distance="300" swimtime="00:03:32.97" />
                    <SPLIT distance="350" swimtime="00:04:09.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" status="DSQ" swimtime="00:05:31.08" resultid="1886" heatid="2405" lane="1" entrytime="00:05:41.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                    <SPLIT distance="100" swimtime="00:01:18.10" />
                    <SPLIT distance="150" swimtime="00:02:04.79" />
                    <SPLIT distance="200" swimtime="00:02:49.96" />
                    <SPLIT distance="250" swimtime="00:03:34.20" />
                    <SPLIT distance="300" swimtime="00:04:17.35" />
                    <SPLIT distance="350" swimtime="00:04:55.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="373" swimtime="00:10:11.57" resultid="1887" heatid="2426" lane="1" entrytime="00:10:02.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.03" />
                    <SPLIT distance="100" swimtime="00:01:11.83" />
                    <SPLIT distance="150" swimtime="00:01:51.25" />
                    <SPLIT distance="200" swimtime="00:02:30.85" />
                    <SPLIT distance="250" swimtime="00:03:10.32" />
                    <SPLIT distance="300" swimtime="00:03:50.11" />
                    <SPLIT distance="350" swimtime="00:04:29.59" />
                    <SPLIT distance="400" swimtime="00:05:08.62" />
                    <SPLIT distance="450" swimtime="00:05:47.67" />
                    <SPLIT distance="500" swimtime="00:06:26.23" />
                    <SPLIT distance="550" swimtime="00:07:04.82" />
                    <SPLIT distance="600" swimtime="00:07:43.39" />
                    <SPLIT distance="650" swimtime="00:08:22.27" />
                    <SPLIT distance="700" swimtime="00:08:59.98" />
                    <SPLIT distance="750" swimtime="00:09:36.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1405" points="406" swimtime="00:02:14.18" resultid="1888" heatid="2414" lane="4" entrytime="00:02:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                    <SPLIT distance="100" swimtime="00:01:03.47" />
                    <SPLIT distance="150" swimtime="00:01:38.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Furuchi Martins" birthdate="2011-10-05" gender="F" nation="BRA" license="367001" athleteid="1962" externalid="367001">
              <RESULTS>
                <RESULT eventid="1087" points="254" swimtime="00:03:12.18" resultid="1963" heatid="2362" lane="4" entrytime="00:03:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.78" />
                    <SPLIT distance="100" swimtime="00:01:39.36" />
                    <SPLIT distance="150" swimtime="00:02:30.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="283" swimtime="00:00:43.18" resultid="1964" heatid="2380" lane="8" entrytime="00:00:41.37" entrycourse="SCM" />
                <RESULT eventid="1232" points="296" swimtime="00:03:21.86" resultid="1965" heatid="2387" lane="1" entrytime="00:03:20.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.04" />
                    <SPLIT distance="150" swimtime="00:02:30.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1444" points="294" swimtime="00:01:33.76" resultid="1966" heatid="2420" lane="6" entrytime="00:01:31.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Biason Santana" birthdate="2009-01-21" gender="M" nation="BRA" license="366969" athleteid="1915" externalid="366969">
              <RESULTS>
                <RESULT eventid="1152" points="374" swimtime="00:02:28.28" resultid="1916" heatid="2374" lane="6" entrytime="00:02:28.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                    <SPLIT distance="100" swimtime="00:01:09.08" />
                    <SPLIT distance="150" swimtime="00:01:45.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1323" points="426" swimtime="00:01:03.48" resultid="1917" heatid="2402" lane="2" entrytime="00:01:02.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="460" swimtime="00:00:28.17" resultid="1918" heatid="2419" lane="3" entrytime="00:00:27.47" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Sol Reolon Gomes" birthdate="2011-02-28" gender="F" nation="BRA" license="392100" athleteid="1951" externalid="392100">
              <RESULTS>
                <RESULT eventid="1113" points="409" swimtime="00:00:34.00" resultid="1952" heatid="2367" lane="8" entrytime="00:00:36.24" entrycourse="SCM" />
                <RESULT comment=" (Horário: 17:36)" eventid="1310" status="DSQ" swimtime="00:01:30.68" resultid="1953" heatid="2399" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="467" swimtime="00:00:29.54" resultid="1954" heatid="2391" lane="3" entrytime="00:00:30.25" entrycourse="SCM" />
                <RESULT eventid="1366" points="357" swimtime="00:01:17.33" resultid="1955" heatid="2409" lane="8" entrytime="00:01:16.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Donato De Morais" birthdate="2009-03-28" gender="F" nation="BRA" license="345588" athleteid="1900" externalid="345588">
              <RESULTS>
                <RESULT eventid="1113" points="356" swimtime="00:00:35.62" resultid="1901" heatid="2367" lane="1" entrytime="00:00:35.40" entrycourse="SCM" />
                <RESULT eventid="1284" points="342" swimtime="00:02:49.93" resultid="1902" heatid="2396" lane="2" entrytime="00:02:41.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.27" />
                    <SPLIT distance="100" swimtime="00:01:23.34" />
                    <SPLIT distance="150" swimtime="00:02:07.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="338" swimtime="00:05:31.86" resultid="1903" heatid="2382" lane="6" entrytime="00:05:28.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                    <SPLIT distance="100" swimtime="00:01:19.11" />
                    <SPLIT distance="150" swimtime="00:02:01.42" />
                    <SPLIT distance="200" swimtime="00:02:44.95" />
                    <SPLIT distance="250" swimtime="00:03:27.91" />
                    <SPLIT distance="300" swimtime="00:04:10.95" />
                    <SPLIT distance="350" swimtime="00:04:53.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="350" swimtime="00:01:17.84" resultid="1904" heatid="2409" lane="7" entrytime="00:01:15.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Schuch Pimpao" birthdate="2010-05-17" gender="M" nation="BRA" license="355586" athleteid="1923" externalid="355586">
              <RESULTS>
                <RESULT eventid="1100" points="352" swimtime="00:00:31.29" resultid="1924" heatid="2365" lane="7" entrytime="00:00:32.47" entrycourse="SCM" />
                <RESULT eventid="1297" points="357" swimtime="00:02:28.81" resultid="1925" heatid="2398" lane="2" entrytime="00:02:30.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                    <SPLIT distance="100" swimtime="00:01:13.24" />
                    <SPLIT distance="150" swimtime="00:01:52.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="358" swimtime="00:01:08.06" resultid="1926" heatid="2410" lane="4" entrytime="00:01:08.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Marques Picolo Vinha" birthdate="2010-07-01" gender="M" nation="BRA" license="366990" athleteid="1967" externalid="366990">
              <RESULTS>
                <RESULT eventid="1219" points="295" swimtime="00:05:18.57" resultid="1968" heatid="2384" lane="3" entrytime="00:05:07.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                    <SPLIT distance="100" swimtime="00:01:11.41" />
                    <SPLIT distance="150" swimtime="00:01:52.44" />
                    <SPLIT distance="200" swimtime="00:02:33.70" />
                    <SPLIT distance="250" swimtime="00:03:15.33" />
                    <SPLIT distance="300" swimtime="00:03:56.61" />
                    <SPLIT distance="350" swimtime="00:04:38.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="276" swimtime="00:11:16.49" resultid="1969" heatid="2425" lane="2" entrytime="00:12:00.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                    <SPLIT distance="100" swimtime="00:01:14.85" />
                    <SPLIT distance="150" swimtime="00:01:57.87" />
                    <SPLIT distance="200" swimtime="00:02:40.82" />
                    <SPLIT distance="250" swimtime="00:03:23.16" />
                    <SPLIT distance="300" swimtime="00:04:06.00" />
                    <SPLIT distance="350" swimtime="00:04:49.70" />
                    <SPLIT distance="400" swimtime="00:05:34.42" />
                    <SPLIT distance="450" swimtime="00:06:18.38" />
                    <SPLIT distance="500" swimtime="00:07:00.63" />
                    <SPLIT distance="550" swimtime="00:07:44.83" />
                    <SPLIT distance="600" swimtime="00:08:27.67" />
                    <SPLIT distance="650" swimtime="00:09:12.06" />
                    <SPLIT distance="700" swimtime="00:09:55.36" />
                    <SPLIT distance="750" swimtime="00:10:37.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Corsine Ferreira" birthdate="2010-03-10" gender="F" nation="BRA" license="353591" athleteid="1939" externalid="353591">
              <RESULTS>
                <RESULT eventid="1113" status="DSQ" swimtime="00:00:35.42" resultid="1940" heatid="2367" lane="2" entrytime="00:00:34.06" entrycourse="SCM" />
                <RESULT eventid="1061" points="316" swimtime="00:22:12.37" resultid="1941" heatid="2358" lane="4" entrytime="00:22:45.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                    <SPLIT distance="100" swimtime="00:01:15.85" />
                    <SPLIT distance="150" swimtime="00:01:56.91" />
                    <SPLIT distance="200" swimtime="00:02:38.43" />
                    <SPLIT distance="250" swimtime="00:03:20.49" />
                    <SPLIT distance="300" swimtime="00:04:03.25" />
                    <SPLIT distance="350" swimtime="00:04:46.36" />
                    <SPLIT distance="400" swimtime="00:05:29.81" />
                    <SPLIT distance="450" swimtime="00:06:13.50" />
                    <SPLIT distance="500" swimtime="00:06:57.35" />
                    <SPLIT distance="550" swimtime="00:07:41.55" />
                    <SPLIT distance="600" swimtime="00:08:25.90" />
                    <SPLIT distance="650" swimtime="00:09:10.88" />
                    <SPLIT distance="700" swimtime="00:09:55.62" />
                    <SPLIT distance="750" swimtime="00:10:40.69" />
                    <SPLIT distance="800" swimtime="00:11:25.65" />
                    <SPLIT distance="850" swimtime="00:12:11.03" />
                    <SPLIT distance="900" swimtime="00:12:56.37" />
                    <SPLIT distance="950" swimtime="00:13:42.02" />
                    <SPLIT distance="1000" swimtime="00:14:27.47" />
                    <SPLIT distance="1050" swimtime="00:15:13.34" />
                    <SPLIT distance="1100" swimtime="00:15:59.39" />
                    <SPLIT distance="1150" swimtime="00:16:45.58" />
                    <SPLIT distance="1200" swimtime="00:17:32.35" />
                    <SPLIT distance="1250" swimtime="00:18:18.95" />
                    <SPLIT distance="1300" swimtime="00:19:05.76" />
                    <SPLIT distance="1350" swimtime="00:19:52.62" />
                    <SPLIT distance="1400" swimtime="00:20:39.16" />
                    <SPLIT distance="1450" swimtime="00:21:25.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="367" swimtime="00:02:46.03" resultid="1942" heatid="2396" lane="6" entrytime="00:02:41.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                    <SPLIT distance="100" swimtime="00:01:19.62" />
                    <SPLIT distance="150" swimtime="00:02:03.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="365" swimtime="00:01:16.76" resultid="1943" heatid="2409" lane="2" entrytime="00:01:14.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Garcia Cavalcante" birthdate="2011-11-21" gender="M" nation="BRA" license="378200" athleteid="1889" externalid="378200">
              <RESULTS>
                <RESULT eventid="1245" points="269" swimtime="00:03:06.11" resultid="1890" heatid="2388" lane="6" entrytime="00:03:10.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.65" />
                    <SPLIT distance="100" swimtime="00:01:28.44" />
                    <SPLIT distance="150" swimtime="00:02:16.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Passafaro" birthdate="2009-02-01" gender="F" nation="BRA" license="370673" athleteid="1905" externalid="370673">
              <RESULTS>
                <RESULT eventid="1139" points="365" swimtime="00:01:10.27" resultid="1906" heatid="2371" lane="5" entrytime="00:01:09.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="278" swimtime="00:01:22.81" resultid="1907" heatid="2400" lane="7" entrytime="00:01:22.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="375" swimtime="00:00:31.79" resultid="1908" heatid="2391" lane="7" entrytime="00:00:30.77" entrycourse="SCM" />
                <RESULT eventid="1418" points="369" swimtime="00:00:33.98" resultid="1909" heatid="2417" lane="6" entrytime="00:00:33.10" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Quental De Meireles" birthdate="2008-11-20" gender="M" nation="BRA" license="392103" athleteid="1956" externalid="392103">
              <RESULTS>
                <RESULT eventid="1271" points="341" swimtime="00:00:28.85" resultid="1957" heatid="2393" lane="2" entrytime="00:00:28.38" entrycourse="SCM" />
                <RESULT eventid="1405" points="398" swimtime="00:02:15.01" resultid="1958" heatid="2415" lane="7" entrytime="00:02:18.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                    <SPLIT distance="100" swimtime="00:01:04.63" />
                    <SPLIT distance="150" swimtime="00:01:40.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="358" swimtime="00:00:30.63" resultid="1959" heatid="2419" lane="1" entrytime="00:00:30.24" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Campelo" birthdate="2011-09-12" gender="M" nation="BRA" license="366963" athleteid="1859" externalid="366963">
              <RESULTS>
                <RESULT eventid="1126" points="440" swimtime="00:00:58.92" resultid="1860" heatid="2370" lane="8" entrytime="00:00:58.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="369" swimtime="00:00:30.81" resultid="1861" heatid="2365" lane="2" entrytime="00:00:31.13" entrycourse="SCM" />
                <RESULT eventid="1297" points="346" swimtime="00:02:30.41" resultid="1862" heatid="2397" lane="5" entrytime="00:02:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="100" swimtime="00:01:11.92" />
                    <SPLIT distance="150" swimtime="00:01:51.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="449" swimtime="00:00:26.31" resultid="1863" heatid="2394" lane="8" entrytime="00:00:26.65" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Chaim" birthdate="2011-05-29" gender="F" nation="BRA" license="370662" athleteid="1933" externalid="370662">
              <RESULTS>
                <RESULT eventid="1139" points="320" swimtime="00:01:13.42" resultid="1934" heatid="2371" lane="6" entrytime="00:01:13.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="288" swimtime="00:05:50.02" resultid="1935" heatid="2382" lane="2" entrytime="00:05:49.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.97" />
                    <SPLIT distance="100" swimtime="00:01:22.27" />
                    <SPLIT distance="150" swimtime="00:02:06.64" />
                    <SPLIT distance="200" swimtime="00:02:51.75" />
                    <SPLIT distance="250" swimtime="00:03:37.53" />
                    <SPLIT distance="300" swimtime="00:04:22.09" />
                    <SPLIT distance="350" swimtime="00:05:06.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="317" swimtime="00:02:41.66" resultid="1936" heatid="2412" lane="6" entrytime="00:02:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                    <SPLIT distance="100" swimtime="00:01:17.28" />
                    <SPLIT distance="150" swimtime="00:02:00.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniela" lastname="Inoue" birthdate="2008-10-31" gender="F" nation="BRA" license="378348" athleteid="1919" externalid="378348">
              <RESULTS>
                <RESULT eventid="1139" points="350" swimtime="00:01:11.27" resultid="1920" heatid="2371" lane="3" entrytime="00:01:10.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="280" swimtime="00:02:48.46" resultid="1921" heatid="2413" lane="1" entrytime="00:02:38.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                    <SPLIT distance="100" swimtime="00:01:19.04" />
                    <SPLIT distance="150" swimtime="00:02:03.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1418" points="287" swimtime="00:00:36.93" resultid="1922" heatid="2416" lane="5" entrytime="00:00:40.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felype" lastname="Gongora Zago" birthdate="2011-09-14" gender="M" nation="BRA" license="392099" athleteid="1949" externalid="392099">
              <RESULTS>
                <RESULT eventid="1379" points="190" swimtime="00:01:23.98" resultid="1950" heatid="2410" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Paiva Boeing" birthdate="2008-01-22" gender="F" nation="BRA" license="318185" athleteid="1891" externalid="318185">
              <RESULTS>
                <RESULT eventid="1191" points="390" swimtime="00:00:38.80" resultid="1892" heatid="2380" lane="7" entrytime="00:00:40.54" entrycourse="SCM" />
                <RESULT eventid="1258" points="407" swimtime="00:00:30.94" resultid="1893" heatid="2391" lane="2" entrytime="00:00:30.71" entrycourse="SCM" />
                <RESULT eventid="1444" points="329" swimtime="00:01:30.26" resultid="1894" heatid="2421" lane="7" entrytime="00:01:24.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietro" lastname="Nabas De Assis" birthdate="2011-07-09" gender="M" nation="BRA" license="366968" athleteid="1927" externalid="366968">
              <RESULTS>
                <RESULT eventid="1178" points="369" swimtime="00:00:34.78" resultid="1928" heatid="2378" lane="1" entrytime="00:00:34.95" entrycourse="SCM" />
                <RESULT eventid="1457" points="384" swimtime="00:01:16.01" resultid="1929" heatid="2423" lane="4" entrytime="00:01:18.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="MARINGÃ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1364" points="576" swimtime="00:03:39.56" resultid="1972" heatid="2407" lane="4" entrytime="00:03:32.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.95" />
                    <SPLIT distance="100" swimtime="00:00:56.33" />
                    <SPLIT distance="150" swimtime="00:01:21.67" />
                    <SPLIT distance="200" swimtime="00:01:48.73" />
                    <SPLIT distance="250" swimtime="00:02:13.95" />
                    <SPLIT distance="300" swimtime="00:02:42.82" />
                    <SPLIT distance="350" swimtime="00:03:09.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1874" number="1" />
                    <RELAYPOSITION athleteid="1864" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1869" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1859" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1485" points="515" swimtime="00:04:08.12" resultid="1973" heatid="2428" lane="4" entrytime="00:03:54.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                    <SPLIT distance="100" swimtime="00:01:07.88" />
                    <SPLIT distance="150" swimtime="00:01:38.56" />
                    <SPLIT distance="200" swimtime="00:02:15.07" />
                    <SPLIT distance="250" swimtime="00:02:42.91" />
                    <SPLIT distance="300" swimtime="00:03:16.04" />
                    <SPLIT distance="350" swimtime="00:03:41.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1874" number="1" />
                    <RELAYPOSITION athleteid="1910" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1869" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1864" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1362" points="440" swimtime="00:04:29.99" resultid="1970" heatid="2406" lane="4" entrytime="00:04:11.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                    <SPLIT distance="100" swimtime="00:01:06.44" />
                    <SPLIT distance="150" swimtime="00:01:37.60" />
                    <SPLIT distance="200" swimtime="00:02:13.01" />
                    <SPLIT distance="250" swimtime="00:02:45.59" />
                    <SPLIT distance="300" swimtime="00:03:23.17" />
                    <SPLIT distance="350" swimtime="00:03:54.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1944" number="1" />
                    <RELAYPOSITION athleteid="1895" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1919" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1951" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1483" points="434" swimtime="00:04:56.25" resultid="1971" heatid="2427" lane="4" entrytime="00:04:44.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                    <SPLIT distance="100" swimtime="00:01:16.63" />
                    <SPLIT distance="150" swimtime="00:01:53.01" />
                    <SPLIT distance="200" swimtime="00:02:35.15" />
                    <SPLIT distance="250" swimtime="00:03:10.36" />
                    <SPLIT distance="300" swimtime="00:03:51.11" />
                    <SPLIT distance="350" swimtime="00:04:22.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1939" number="1" />
                    <RELAYPOSITION athleteid="1895" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1944" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1951" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="MARINGÃÂ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1204" status="DSQ" swimtime="00:02:00.68" resultid="1974" heatid="2381" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.78" />
                    <SPLIT distance="100" swimtime="00:01:05.47" />
                    <SPLIT distance="150" swimtime="00:01:31.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1939" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="1910" number="2" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION athleteid="1864" number="3" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION athleteid="1895" number="4" reactiontime="0" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="689" nation="BRA" region="PR" clubid="1512" name="Seleção De Cascavel/PR" shortname="Cascavel">
          <ATHLETES>
            <ATHLETE firstname="Giovanna" lastname="Bertelli Weirich" birthdate="2011-03-18" gender="F" nation="BRA" license="369534" athleteid="1564" externalid="369534">
              <RESULTS>
                <RESULT eventid="1165" points="407" swimtime="00:02:41.31" resultid="1565" heatid="2376" lane="6" entrytime="00:02:51.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                    <SPLIT distance="100" swimtime="00:01:16.30" />
                    <SPLIT distance="150" swimtime="00:01:58.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="470" swimtime="00:04:57.48" resultid="1566" heatid="2383" lane="6" entrytime="00:05:01.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="100" swimtime="00:01:10.64" />
                    <SPLIT distance="150" swimtime="00:01:48.49" />
                    <SPLIT distance="200" swimtime="00:02:26.58" />
                    <SPLIT distance="250" swimtime="00:03:04.29" />
                    <SPLIT distance="300" swimtime="00:03:42.64" />
                    <SPLIT distance="350" swimtime="00:04:20.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="428" swimtime="00:05:43.38" resultid="1567" heatid="2403" lane="2" entrytime="00:06:03.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                    <SPLIT distance="100" swimtime="00:01:18.81" />
                    <SPLIT distance="150" swimtime="00:02:03.00" />
                    <SPLIT distance="200" swimtime="00:02:46.37" />
                    <SPLIT distance="250" swimtime="00:03:34.75" />
                    <SPLIT distance="300" swimtime="00:04:25.03" />
                    <SPLIT distance="350" swimtime="00:05:05.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1418" points="365" swimtime="00:00:34.11" resultid="1568" heatid="2417" lane="8" entrytime="00:00:35.05" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Gamero Prado" birthdate="2007-05-16" gender="F" nation="BRA" license="305973" athleteid="1513" externalid="305973">
              <RESULTS>
                <RESULT eventid="1165" points="360" swimtime="00:02:48.03" resultid="1514" heatid="2376" lane="3" entrytime="00:02:49.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                    <SPLIT distance="100" swimtime="00:01:17.49" />
                    <SPLIT distance="150" swimtime="00:02:01.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1061" points="323" swimtime="00:22:03.35" resultid="1515" heatid="2359" lane="3" entrytime="00:20:28.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                    <SPLIT distance="100" swimtime="00:01:12.54" />
                    <SPLIT distance="150" swimtime="00:01:51.19" />
                    <SPLIT distance="200" swimtime="00:02:30.31" />
                    <SPLIT distance="250" swimtime="00:03:11.03" />
                    <SPLIT distance="300" swimtime="00:03:53.58" />
                    <SPLIT distance="350" swimtime="00:04:36.32" />
                    <SPLIT distance="400" swimtime="00:05:18.37" />
                    <SPLIT distance="450" swimtime="00:06:00.38" />
                    <SPLIT distance="500" swimtime="00:06:43.37" />
                    <SPLIT distance="550" swimtime="00:07:24.93" />
                    <SPLIT distance="600" swimtime="00:08:06.85" />
                    <SPLIT distance="650" swimtime="00:08:49.56" />
                    <SPLIT distance="700" swimtime="00:09:32.15" />
                    <SPLIT distance="750" swimtime="00:10:15.21" />
                    <SPLIT distance="800" swimtime="00:10:58.71" />
                    <SPLIT distance="850" swimtime="00:11:40.70" />
                    <SPLIT distance="900" swimtime="00:12:23.58" />
                    <SPLIT distance="950" swimtime="00:13:06.41" />
                    <SPLIT distance="1000" swimtime="00:13:49.14" />
                    <SPLIT distance="1050" swimtime="00:14:32.53" />
                    <SPLIT distance="1100" swimtime="00:15:16.58" />
                    <SPLIT distance="1150" swimtime="00:15:59.89" />
                    <SPLIT distance="1200" swimtime="00:16:43.29" />
                    <SPLIT distance="1250" swimtime="00:17:27.32" />
                    <SPLIT distance="1300" swimtime="00:18:10.14" />
                    <SPLIT distance="1350" swimtime="00:18:53.20" />
                    <SPLIT distance="1400" swimtime="00:19:35.86" />
                    <SPLIT distance="1450" swimtime="00:20:18.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="390" swimtime="00:01:13.93" resultid="1516" heatid="2400" lane="3" entrytime="00:01:14.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1418" points="375" swimtime="00:00:33.80" resultid="1517" heatid="2417" lane="2" entrytime="00:00:33.54" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Assakura" birthdate="2010-06-29" gender="F" nation="BRA" license="376473" athleteid="1592" externalid="376473">
              <RESULTS>
                <RESULT eventid="1087" points="449" swimtime="00:02:39.04" resultid="1593" heatid="2363" lane="6" entrytime="00:02:42.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.69" />
                    <SPLIT distance="100" swimtime="00:01:17.24" />
                    <SPLIT distance="150" swimtime="00:02:01.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="385" swimtime="00:00:38.99" resultid="1594" heatid="2380" lane="2" entrytime="00:00:40.33" entrycourse="SCM" />
                <RESULT eventid="1232" points="505" swimtime="00:02:48.96" resultid="1595" heatid="2387" lane="5" entrytime="00:02:57.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.73" />
                    <SPLIT distance="100" swimtime="00:01:21.16" />
                    <SPLIT distance="150" swimtime="00:02:04.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1444" points="388" swimtime="00:01:25.46" resultid="1596" heatid="2421" lane="2" entrytime="00:01:24.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Rinaldini" birthdate="2009-04-09" gender="M" nation="BRA" license="348289" athleteid="1523" externalid="348289">
              <RESULTS>
                <RESULT eventid="1152" points="526" swimtime="00:02:12.30" resultid="1524" heatid="2374" lane="4" entrytime="00:02:15.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                    <SPLIT distance="100" swimtime="00:01:03.14" />
                    <SPLIT distance="150" swimtime="00:01:37.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="588" swimtime="00:04:13.21" resultid="1525" heatid="2385" lane="3" entrytime="00:04:18.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                    <SPLIT distance="100" swimtime="00:01:00.82" />
                    <SPLIT distance="150" swimtime="00:01:32.85" />
                    <SPLIT distance="200" swimtime="00:02:05.57" />
                    <SPLIT distance="250" swimtime="00:02:37.81" />
                    <SPLIT distance="300" swimtime="00:03:10.18" />
                    <SPLIT distance="350" swimtime="00:03:42.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="537" swimtime="00:04:48.71" resultid="1526" heatid="2405" lane="5" entrytime="00:04:56.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                    <SPLIT distance="100" swimtime="00:01:04.22" />
                    <SPLIT distance="150" swimtime="00:01:42.40" />
                    <SPLIT distance="200" swimtime="00:02:20.12" />
                    <SPLIT distance="250" swimtime="00:03:01.41" />
                    <SPLIT distance="300" swimtime="00:03:43.88" />
                    <SPLIT distance="350" swimtime="00:04:16.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="577" swimtime="00:08:48.90" resultid="1527" heatid="2426" lane="3" entrytime="00:08:55.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                    <SPLIT distance="100" swimtime="00:01:02.64" />
                    <SPLIT distance="150" swimtime="00:01:35.41" />
                    <SPLIT distance="200" swimtime="00:02:09.00" />
                    <SPLIT distance="250" swimtime="00:02:42.53" />
                    <SPLIT distance="300" swimtime="00:03:16.31" />
                    <SPLIT distance="350" swimtime="00:03:49.61" />
                    <SPLIT distance="400" swimtime="00:04:22.90" />
                    <SPLIT distance="450" swimtime="00:04:55.99" />
                    <SPLIT distance="500" swimtime="00:05:29.19" />
                    <SPLIT distance="550" swimtime="00:06:02.74" />
                    <SPLIT distance="600" swimtime="00:06:36.70" />
                    <SPLIT distance="650" swimtime="00:07:10.15" />
                    <SPLIT distance="700" swimtime="00:07:43.86" />
                    <SPLIT distance="750" swimtime="00:08:16.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luann" lastname="Miguel Mazur" birthdate="2007-01-10" gender="M" nation="BRA" license="365682" athleteid="1546" externalid="365682">
              <RESULTS>
                <RESULT eventid="1178" points="397" swimtime="00:00:33.93" resultid="1547" heatid="2378" lane="6" entrytime="00:00:33.46" entrycourse="SCM" />
                <RESULT eventid="1349" points="487" swimtime="00:04:58.43" resultid="1548" heatid="2405" lane="3" entrytime="00:04:57.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                    <SPLIT distance="100" swimtime="00:01:07.83" />
                    <SPLIT distance="150" swimtime="00:01:45.93" />
                    <SPLIT distance="200" swimtime="00:02:23.22" />
                    <SPLIT distance="250" swimtime="00:03:04.77" />
                    <SPLIT distance="300" swimtime="00:03:47.09" />
                    <SPLIT distance="350" swimtime="00:04:22.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="451" swimtime="00:01:12.07" resultid="1549" heatid="2424" lane="6" entrytime="00:01:10.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Alves Serafini" birthdate="2008-04-15" gender="M" nation="BRA" license="351644" athleteid="1601" externalid="351644">
              <RESULTS>
                <RESULT eventid="1152" points="503" swimtime="00:02:14.29" resultid="1602" heatid="2374" lane="5" entrytime="00:02:21.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.15" />
                    <SPLIT distance="100" swimtime="00:01:02.97" />
                    <SPLIT distance="150" swimtime="00:01:36.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1323" points="482" swimtime="00:01:00.90" resultid="1603" heatid="2402" lane="3" entrytime="00:01:01.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="422" swimtime="00:00:28.99" resultid="1604" heatid="2418" lane="6" entrytime="00:00:36.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Sehn Uren" birthdate="2009-10-15" gender="F" nation="BRA" license="357159" athleteid="1533" externalid="357159">
              <RESULTS>
                <RESULT eventid="1139" points="409" swimtime="00:01:07.68" resultid="1534" heatid="2372" lane="8" entrytime="00:01:08.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="432" swimtime="00:02:37.30" resultid="1535" heatid="2396" lane="3" entrytime="00:02:40.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.41" />
                    <SPLIT distance="100" swimtime="00:01:18.06" />
                    <SPLIT distance="150" swimtime="00:01:57.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="424" swimtime="00:05:44.54" resultid="1536" heatid="2403" lane="6" entrytime="00:05:57.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.98" />
                    <SPLIT distance="100" swimtime="00:01:22.53" />
                    <SPLIT distance="150" swimtime="00:02:08.73" />
                    <SPLIT distance="200" swimtime="00:02:51.61" />
                    <SPLIT distance="250" swimtime="00:03:38.59" />
                    <SPLIT distance="300" swimtime="00:04:25.98" />
                    <SPLIT distance="350" swimtime="00:05:06.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="360" swimtime="00:01:17.10" resultid="1537" heatid="2408" lane="4" entrytime="00:01:16.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Breno" lastname="Zanella Janke" birthdate="2011-04-26" gender="M" nation="BRA" license="365697" athleteid="1559" externalid="365697">
              <RESULTS>
                <RESULT eventid="1074" points="414" swimtime="00:02:27.00" resultid="1560" heatid="2361" lane="8" entrytime="00:02:28.15" entrycourse="SCM" />
                <RESULT eventid="1178" points="350" swimtime="00:00:35.39" resultid="1561" heatid="2378" lane="8" entrytime="00:00:35.63" entrycourse="SCM" />
                <RESULT eventid="1271" points="390" swimtime="00:00:27.57" resultid="1562" heatid="2392" lane="4" entrytime="00:00:30.00" entrycourse="SCM" />
                <RESULT eventid="1405" points="397" swimtime="00:02:15.18" resultid="1563" heatid="2414" lane="3" entrytime="00:02:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.70" />
                    <SPLIT distance="100" swimtime="00:01:03.45" />
                    <SPLIT distance="150" swimtime="00:01:39.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raul" lastname="Bonamigo" birthdate="2010-12-01" gender="M" nation="BRA" license="344397" athleteid="1597" externalid="344397">
              <RESULTS>
                <RESULT eventid="1100" points="361" swimtime="00:00:31.05" resultid="1598" heatid="2364" lane="4" entrytime="00:00:35.00" entrycourse="SCM" />
                <RESULT eventid="1297" points="384" swimtime="00:02:25.32" resultid="1599" heatid="2398" lane="6" entrytime="00:02:27.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.01" />
                    <SPLIT distance="100" swimtime="00:01:10.61" />
                    <SPLIT distance="150" swimtime="00:01:48.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="369" swimtime="00:01:07.35" resultid="1600" heatid="2411" lane="1" entrytime="00:01:07.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hendrik" lastname="Alteiro Groenwold" birthdate="2011-03-23" gender="M" nation="BRA" license="365756" athleteid="1550" externalid="365756">
              <RESULTS>
                <RESULT eventid="1152" points="425" swimtime="00:02:22.02" resultid="1551" heatid="2374" lane="2" entrytime="00:02:42.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                    <SPLIT distance="100" swimtime="00:01:07.16" />
                    <SPLIT distance="150" swimtime="00:01:44.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1323" points="386" swimtime="00:01:05.58" resultid="1552" heatid="2402" lane="8" entrytime="00:01:05.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1405" points="446" swimtime="00:02:09.99" resultid="1553" heatid="2415" lane="2" entrytime="00:02:11.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                    <SPLIT distance="100" swimtime="00:01:02.32" />
                    <SPLIT distance="150" swimtime="00:01:35.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emanuel" lastname="Ranieri" birthdate="2011-01-24" gender="M" nation="BRA" license="390838" athleteid="1605" externalid="390838">
              <RESULTS>
                <RESULT eventid="1126" points="353" swimtime="00:01:03.41" resultid="1606" heatid="2369" lane="7" entrytime="00:01:04.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="298" swimtime="00:02:38.09" resultid="1607" heatid="2398" lane="1" entrytime="00:02:40.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                    <SPLIT distance="100" swimtime="00:01:18.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="277" swimtime="00:01:14.09" resultid="1608" heatid="2410" lane="3" entrytime="00:01:14.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juan" lastname="Balduíno" birthdate="2009-06-24" gender="M" nation="BRA" license="370764" athleteid="1578" externalid="370764">
              <RESULTS>
                <RESULT eventid="1100" points="398" swimtime="00:00:30.05" resultid="1579" heatid="2365" lane="6" entrytime="00:00:30.91" entrycourse="SCM" />
                <RESULT eventid="1323" points="472" swimtime="00:01:01.35" resultid="1580" heatid="2402" lane="7" entrytime="00:01:02.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="408" swimtime="00:01:05.15" resultid="1581" heatid="2411" lane="2" entrytime="00:01:06.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Tolentino Smarczewski" birthdate="2008-09-01" gender="M" nation="BRA" license="378818" athleteid="1582" externalid="378818">
              <RESULTS>
                <RESULT eventid="1245" points="415" swimtime="00:02:41.09" resultid="1583" heatid="2389" lane="1" entrytime="00:02:41.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                    <SPLIT distance="100" swimtime="00:01:18.33" />
                    <SPLIT distance="150" swimtime="00:01:59.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" status="DSQ" swimtime="00:00:28.50" resultid="1584" heatid="2393" lane="3" entrytime="00:00:28.14" entrycourse="SCM" />
                <RESULT eventid="1457" points="335" swimtime="00:01:19.55" resultid="1585" heatid="2424" lane="8" entrytime="00:01:15.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1405" points="481" swimtime="00:02:06.75" resultid="1586" heatid="2415" lane="6" entrytime="00:02:09.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.87" />
                    <SPLIT distance="100" swimtime="00:01:01.70" />
                    <SPLIT distance="150" swimtime="00:01:34.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amanda" lastname="Borille Busetti" birthdate="2010-02-17" gender="F" nation="BRA" license="392830" athleteid="1618" externalid="392830">
              <RESULTS>
                <RESULT eventid="1139" points="417" swimtime="00:01:07.23" resultid="1619" heatid="2371" lane="4" entrytime="00:01:08.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="389" swimtime="00:00:31.39" resultid="1620" heatid="2391" lane="8" entrytime="00:00:31.52" entrycourse="SCM" />
                <RESULT eventid="1366" points="307" swimtime="00:01:21.34" resultid="1621" heatid="2408" lane="7" entrytime="00:01:23.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="357" swimtime="00:02:35.36" resultid="1622" heatid="2413" lane="2" entrytime="00:02:32.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                    <SPLIT distance="100" swimtime="00:01:15.97" />
                    <SPLIT distance="150" swimtime="00:01:56.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Colaco Da Conceicao" birthdate="2011-05-25" gender="F" nation="BRA" license="369535" athleteid="1569" externalid="369535">
              <RESULTS>
                <RESULT eventid="1139" points="357" swimtime="00:01:10.83" resultid="1570" heatid="2372" lane="1" entrytime="00:01:08.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1061" points="347" swimtime="00:21:32.44" resultid="1571" heatid="2359" lane="7" entrytime="00:21:45.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:30.63" />
                    <SPLIT distance="100" swimtime="00:03:09.78" />
                    <SPLIT distance="150" swimtime="00:03:49.20" />
                    <SPLIT distance="200" swimtime="00:04:29.15" />
                    <SPLIT distance="250" swimtime="00:05:08.92" />
                    <SPLIT distance="300" swimtime="00:05:48.15" />
                    <SPLIT distance="350" swimtime="00:06:28.83" />
                    <SPLIT distance="400" swimtime="00:07:09.17" />
                    <SPLIT distance="450" swimtime="00:07:50.29" />
                    <SPLIT distance="500" swimtime="00:08:31.54" />
                    <SPLIT distance="550" swimtime="00:09:12.39" />
                    <SPLIT distance="600" swimtime="00:09:53.89" />
                    <SPLIT distance="650" swimtime="00:10:35.31" />
                    <SPLIT distance="700" swimtime="00:11:16.84" />
                    <SPLIT distance="750" swimtime="00:11:58.03" />
                    <SPLIT distance="800" swimtime="00:12:39.22" />
                    <SPLIT distance="850" swimtime="00:13:21.30" />
                    <SPLIT distance="900" swimtime="00:14:02.63" />
                    <SPLIT distance="950" swimtime="00:14:44.09" />
                    <SPLIT distance="1000" swimtime="00:15:25.42" />
                    <SPLIT distance="1050" swimtime="00:16:06.90" />
                    <SPLIT distance="1100" swimtime="00:16:48.73" />
                    <SPLIT distance="1150" swimtime="00:17:30.97" />
                    <SPLIT distance="1200" swimtime="00:18:12.24" />
                    <SPLIT distance="1250" swimtime="00:18:53.30" />
                    <SPLIT distance="1300" swimtime="00:19:33.49" />
                    <SPLIT distance="1350" swimtime="00:20:15.67" />
                    <SPLIT distance="1400" swimtime="00:20:55.14" />
                    <SPLIT distance="1450" swimtime="00:21:32.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="403" swimtime="00:05:12.90" resultid="1572" heatid="2383" lane="3" entrytime="00:04:57.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                    <SPLIT distance="100" swimtime="00:01:11.84" />
                    <SPLIT distance="150" swimtime="00:01:51.23" />
                    <SPLIT distance="200" swimtime="00:02:30.81" />
                    <SPLIT distance="250" swimtime="00:03:11.46" />
                    <SPLIT distance="300" swimtime="00:03:52.62" />
                    <SPLIT distance="350" swimtime="00:04:32.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="384" swimtime="00:02:31.64" resultid="1573" heatid="2413" lane="7" entrytime="00:02:33.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                    <SPLIT distance="100" swimtime="00:01:12.13" />
                    <SPLIT distance="150" swimtime="00:01:52.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Stein Duarte" birthdate="2010-10-03" gender="F" nation="BRA" license="351635" athleteid="1528" externalid="351635">
              <RESULTS>
                <RESULT eventid="1087" points="470" swimtime="00:02:36.70" resultid="1529" heatid="2363" lane="5" entrytime="00:02:37.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                    <SPLIT distance="100" swimtime="00:01:12.15" />
                    <SPLIT distance="150" swimtime="00:01:58.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="440" swimtime="00:00:33.19" resultid="1530" heatid="2367" lane="3" entrytime="00:00:33.48" entrycourse="SCM" />
                <RESULT eventid="1284" points="450" swimtime="00:02:35.11" resultid="1531" heatid="2396" lane="5" entrytime="00:02:36.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                    <SPLIT distance="100" swimtime="00:01:15.92" />
                    <SPLIT distance="150" swimtime="00:01:56.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="452" swimtime="00:01:11.48" resultid="1532" heatid="2409" lane="5" entrytime="00:01:10.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Zimmermann" birthdate="2010-01-19" gender="M" nation="BRA" license="357160" athleteid="1538" externalid="357160">
              <RESULTS>
                <RESULT eventid="1074" points="507" swimtime="00:02:17.47" resultid="1539" heatid="2361" lane="3" entrytime="00:02:20.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.69" />
                    <SPLIT distance="100" swimtime="00:01:46.36" />
                    <SPLIT distance="150" swimtime="00:02:17.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="471" swimtime="00:02:15.71" resultid="1540" heatid="2398" lane="5" entrytime="00:02:19.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                    <SPLIT distance="100" swimtime="00:01:06.17" />
                    <SPLIT distance="150" swimtime="00:01:41.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="522" swimtime="00:09:06.91" resultid="1541" heatid="2426" lane="5" entrytime="00:08:53.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.62" />
                    <SPLIT distance="100" swimtime="00:01:02.04" />
                    <SPLIT distance="150" swimtime="00:01:36.16" />
                    <SPLIT distance="200" swimtime="00:02:10.73" />
                    <SPLIT distance="250" swimtime="00:02:45.35" />
                    <SPLIT distance="300" swimtime="00:03:20.05" />
                    <SPLIT distance="350" swimtime="00:03:54.82" />
                    <SPLIT distance="400" swimtime="00:04:29.80" />
                    <SPLIT distance="450" swimtime="00:05:04.73" />
                    <SPLIT distance="500" swimtime="00:05:39.74" />
                    <SPLIT distance="550" swimtime="00:06:14.40" />
                    <SPLIT distance="600" swimtime="00:06:49.86" />
                    <SPLIT distance="650" swimtime="00:07:24.42" />
                    <SPLIT distance="700" swimtime="00:07:58.93" />
                    <SPLIT distance="750" swimtime="00:08:32.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Do Prado Martins" birthdate="2008-10-17" gender="F" nation="BRA" license="369419" athleteid="1554" externalid="369419">
              <RESULTS>
                <RESULT eventid="1087" points="502" swimtime="00:02:33.25" resultid="1555" heatid="2363" lane="4" entrytime="00:02:37.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                    <SPLIT distance="100" swimtime="00:01:12.37" />
                    <SPLIT distance="150" swimtime="00:01:55.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="501" swimtime="00:02:49.40" resultid="1556" heatid="2387" lane="4" entrytime="00:02:54.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                    <SPLIT distance="100" swimtime="00:01:20.77" />
                    <SPLIT distance="150" swimtime="00:02:04.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="479" swimtime="00:05:30.78" resultid="1557" heatid="2403" lane="5" entrytime="00:05:33.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.35" />
                    <SPLIT distance="100" swimtime="00:01:14.85" />
                    <SPLIT distance="150" swimtime="00:01:58.34" />
                    <SPLIT distance="200" swimtime="00:02:40.80" />
                    <SPLIT distance="250" swimtime="00:03:25.87" />
                    <SPLIT distance="300" swimtime="00:04:12.54" />
                    <SPLIT distance="350" swimtime="00:04:52.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1444" points="484" swimtime="00:01:19.40" resultid="1558" heatid="2421" lane="4" entrytime="00:01:19.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Claudio" lastname="Rohnelt" birthdate="2010-03-08" gender="M" nation="BRA" license="357954" athleteid="1542" externalid="357954">
              <RESULTS>
                <RESULT eventid="1126" points="387" swimtime="00:01:01.52" resultid="1543" heatid="2369" lane="6" entrytime="00:01:03.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="428" swimtime="00:04:41.46" resultid="1544" heatid="2384" lane="5" entrytime="00:04:59.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                    <SPLIT distance="100" swimtime="00:01:07.59" />
                    <SPLIT distance="150" swimtime="00:01:43.50" />
                    <SPLIT distance="200" swimtime="00:02:19.31" />
                    <SPLIT distance="250" swimtime="00:02:55.32" />
                    <SPLIT distance="300" swimtime="00:03:31.61" />
                    <SPLIT distance="350" swimtime="00:04:07.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="315" swimtime="00:00:31.95" resultid="1545" heatid="2418" lane="5" entrytime="00:00:33.63" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Flavia" lastname="De Metz" birthdate="2011-01-07" gender="F" nation="BRA" license="390846" athleteid="1609" externalid="390846">
              <RESULTS>
                <RESULT eventid="1061" points="310" swimtime="00:22:21.03" resultid="1610" heatid="2359" lane="2" entrytime="00:21:42.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                    <SPLIT distance="100" swimtime="00:01:13.41" />
                    <SPLIT distance="150" swimtime="00:01:52.51" />
                    <SPLIT distance="200" swimtime="00:02:32.61" />
                    <SPLIT distance="250" swimtime="00:03:13.96" />
                    <SPLIT distance="300" swimtime="00:03:55.59" />
                    <SPLIT distance="350" swimtime="00:04:38.13" />
                    <SPLIT distance="400" swimtime="00:05:19.79" />
                    <SPLIT distance="450" swimtime="00:06:02.11" />
                    <SPLIT distance="500" swimtime="00:06:43.78" />
                    <SPLIT distance="550" swimtime="00:07:26.31" />
                    <SPLIT distance="600" swimtime="00:08:08.69" />
                    <SPLIT distance="650" swimtime="00:08:50.83" />
                    <SPLIT distance="700" swimtime="00:09:34.14" />
                    <SPLIT distance="750" swimtime="00:10:18.02" />
                    <SPLIT distance="800" swimtime="00:11:01.19" />
                    <SPLIT distance="850" swimtime="00:11:45.19" />
                    <SPLIT distance="900" swimtime="00:12:28.66" />
                    <SPLIT distance="950" swimtime="00:13:13.07" />
                    <SPLIT distance="1000" swimtime="00:13:56.79" />
                    <SPLIT distance="1050" swimtime="00:14:41.21" />
                    <SPLIT distance="1100" swimtime="00:15:25.38" />
                    <SPLIT distance="1150" swimtime="00:16:08.65" />
                    <SPLIT distance="1200" swimtime="00:16:53.24" />
                    <SPLIT distance="1250" swimtime="00:17:37.50" />
                    <SPLIT distance="1300" swimtime="00:18:21.15" />
                    <SPLIT distance="1350" swimtime="00:19:03.69" />
                    <SPLIT distance="1400" swimtime="00:19:47.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="349" swimtime="00:02:48.86" resultid="1611" heatid="2396" lane="7" entrytime="00:02:44.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                    <SPLIT distance="100" swimtime="00:01:21.78" />
                    <SPLIT distance="150" swimtime="00:02:05.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="419" swimtime="00:05:08.93" resultid="1612" heatid="2382" lane="4" entrytime="00:05:12.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                    <SPLIT distance="100" swimtime="00:01:11.63" />
                    <SPLIT distance="150" swimtime="00:01:50.63" />
                    <SPLIT distance="200" swimtime="00:02:30.05" />
                    <SPLIT distance="250" swimtime="00:03:09.71" />
                    <SPLIT distance="300" swimtime="00:03:50.05" />
                    <SPLIT distance="350" swimtime="00:04:29.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="452" swimtime="00:02:23.65" resultid="1613" heatid="2413" lane="3" entrytime="00:02:24.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                    <SPLIT distance="100" swimtime="00:01:08.78" />
                    <SPLIT distance="150" swimtime="00:01:46.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Mariotti De Castro" birthdate="2008-06-27" gender="M" nation="BRA" license="329200" athleteid="1518" externalid="329200">
              <RESULTS>
                <RESULT eventid="1074" points="575" swimtime="00:02:11.82" resultid="1519" heatid="2361" lane="5" entrytime="00:02:16.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.43" />
                    <SPLIT distance="100" swimtime="00:01:02.03" />
                    <SPLIT distance="150" swimtime="00:01:41.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="632" swimtime="00:04:07.26" resultid="1520" heatid="2385" lane="4" entrytime="00:04:03.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.34" />
                    <SPLIT distance="100" swimtime="00:00:58.80" />
                    <SPLIT distance="150" swimtime="00:01:29.88" />
                    <SPLIT distance="200" swimtime="00:02:01.73" />
                    <SPLIT distance="250" swimtime="00:02:32.65" />
                    <SPLIT distance="300" swimtime="00:03:03.53" />
                    <SPLIT distance="350" swimtime="00:03:35.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="619" swimtime="00:04:35.50" resultid="1521" heatid="2405" lane="4" entrytime="00:04:36.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.21" />
                    <SPLIT distance="100" swimtime="00:01:01.70" />
                    <SPLIT distance="150" swimtime="00:01:37.31" />
                    <SPLIT distance="200" swimtime="00:02:12.61" />
                    <SPLIT distance="250" swimtime="00:02:52.53" />
                    <SPLIT distance="300" swimtime="00:03:32.95" />
                    <SPLIT distance="350" swimtime="00:04:05.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="644" swimtime="00:08:29.92" resultid="1522" heatid="2426" lane="4" entrytime="00:08:38.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.89" />
                    <SPLIT distance="100" swimtime="00:01:00.05" />
                    <SPLIT distance="150" swimtime="00:01:32.15" />
                    <SPLIT distance="200" swimtime="00:02:04.99" />
                    <SPLIT distance="250" swimtime="00:02:37.29" />
                    <SPLIT distance="300" swimtime="00:03:09.60" />
                    <SPLIT distance="350" swimtime="00:03:42.24" />
                    <SPLIT distance="400" swimtime="00:04:15.01" />
                    <SPLIT distance="450" swimtime="00:04:46.80" />
                    <SPLIT distance="500" swimtime="00:05:18.68" />
                    <SPLIT distance="550" swimtime="00:05:50.44" />
                    <SPLIT distance="600" swimtime="00:06:22.94" />
                    <SPLIT distance="650" swimtime="00:06:55.11" />
                    <SPLIT distance="700" swimtime="00:07:28.03" />
                    <SPLIT distance="750" swimtime="00:07:59.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Danilo" lastname="Rodrigues" birthdate="2011-05-23" gender="M" nation="BRA" license="370763" athleteid="1574" externalid="370763">
              <RESULTS>
                <RESULT eventid="1126" points="338" swimtime="00:01:04.34" resultid="1575" heatid="2368" lane="5" entrytime="00:01:07.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1245" points="325" swimtime="00:02:54.64" resultid="1576" heatid="2389" lane="8" entrytime="00:03:01.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.29" />
                    <SPLIT distance="100" swimtime="00:01:24.94" />
                    <SPLIT distance="150" swimtime="00:02:10.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="279" swimtime="00:00:33.27" resultid="1577" heatid="2418" lane="3" entrytime="00:00:33.63" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Luisa Lottermann" birthdate="2011-08-26" gender="F" nation="BRA" license="382238" athleteid="1587" externalid="382238">
              <RESULTS>
                <RESULT eventid="1165" points="258" swimtime="00:03:07.66" resultid="1588" heatid="2376" lane="7" entrytime="00:03:07.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.93" />
                    <SPLIT distance="100" swimtime="00:01:30.92" />
                    <SPLIT distance="150" swimtime="00:02:19.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="333" swimtime="00:00:40.90" resultid="1589" heatid="2379" lane="4" entrytime="00:00:41.83" entrycourse="SCM" />
                <RESULT eventid="1232" points="421" swimtime="00:02:59.47" resultid="1590" heatid="2387" lane="6" entrytime="00:03:03.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.91" />
                    <SPLIT distance="100" swimtime="00:01:27.62" />
                    <SPLIT distance="150" swimtime="00:02:13.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1444" points="345" swimtime="00:01:28.83" resultid="1591" heatid="2420" lane="5" entrytime="00:01:28.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Ramirez Vasconcelos" birthdate="2011-04-06" gender="M" nation="BRA" license="392013" athleteid="1614" externalid="392013">
              <RESULTS>
                <RESULT eventid="1178" points="332" swimtime="00:00:36.03" resultid="1615" heatid="2377" lane="5" entrytime="00:00:37.99" entrycourse="SCM" />
                <RESULT eventid="1245" points="355" swimtime="00:02:49.61" resultid="1616" heatid="2388" lane="5" entrytime="00:03:08.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                    <SPLIT distance="100" swimtime="00:01:20.22" />
                    <SPLIT distance="150" swimtime="00:02:04.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="384" swimtime="00:01:16.03" resultid="1617" heatid="2423" lane="3" entrytime="00:01:21.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1364" points="541" swimtime="00:03:44.28" resultid="1625" heatid="2407" lane="6" entrytime="00:03:49.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.66" />
                    <SPLIT distance="100" swimtime="00:00:54.87" />
                    <SPLIT distance="150" swimtime="00:01:22.24" />
                    <SPLIT distance="200" swimtime="00:01:52.23" />
                    <SPLIT distance="250" swimtime="00:02:19.11" />
                    <SPLIT distance="300" swimtime="00:02:48.03" />
                    <SPLIT distance="350" swimtime="00:03:14.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1518" number="1" />
                    <RELAYPOSITION athleteid="1601" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1538" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1578" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1485" points="503" swimtime="00:04:10.17" resultid="1626" heatid="2428" lane="6" entrytime="00:04:23.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                    <SPLIT distance="100" swimtime="00:01:03.30" />
                    <SPLIT distance="150" swimtime="00:01:37.55" />
                    <SPLIT distance="200" swimtime="00:02:15.23" />
                    <SPLIT distance="250" swimtime="00:02:43.76" />
                    <SPLIT distance="300" swimtime="00:03:15.89" />
                    <SPLIT distance="350" swimtime="00:03:42.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1538" number="1" />
                    <RELAYPOSITION athleteid="1546" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1601" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1518" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1362" points="475" swimtime="00:04:23.28" resultid="1623" heatid="2406" lane="6" entrytime="00:04:39.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                    <SPLIT distance="100" swimtime="00:01:06.68" />
                    <SPLIT distance="150" swimtime="00:01:36.81" />
                    <SPLIT distance="200" swimtime="00:02:10.15" />
                    <SPLIT distance="250" swimtime="00:02:42.64" />
                    <SPLIT distance="300" swimtime="00:03:18.43" />
                    <SPLIT distance="350" swimtime="00:03:49.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1528" number="1" />
                    <RELAYPOSITION athleteid="1592" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1513" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1554" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1483" points="451" swimtime="00:04:52.35" resultid="1624" heatid="2427" lane="3" entrytime="00:05:08.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                    <SPLIT distance="100" swimtime="00:01:12.54" />
                    <SPLIT distance="150" swimtime="00:01:49.47" />
                    <SPLIT distance="200" swimtime="00:02:32.25" />
                    <SPLIT distance="250" swimtime="00:03:06.08" />
                    <SPLIT distance="300" swimtime="00:03:46.64" />
                    <SPLIT distance="350" swimtime="00:04:18.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1528" number="1" />
                    <RELAYPOSITION athleteid="1554" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1513" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1592" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1204" points="450" swimtime="00:02:04.11" resultid="1627" heatid="2381" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                    <SPLIT distance="100" swimtime="00:01:09.99" />
                    <SPLIT distance="150" swimtime="00:01:38.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1528" number="1" />
                    <RELAYPOSITION athleteid="1554" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1601" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1518" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="1485" nation="BRA" region="PR" clubid="1487" name="Seleção De Campo Mourão/PR" shortname="Campo Mourão">
          <ATHLETES>
            <ATHLETE firstname="Kenzo" lastname="Kimura" birthdate="2010-04-23" gender="M" nation="BRA" license="403429" athleteid="1504" externalid="403429">
              <RESULTS>
                <RESULT eventid="1126" points="235" swimtime="00:01:12.65" resultid="1505" heatid="2368" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="235" swimtime="00:00:32.65" resultid="1506" heatid="2392" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Gabrieli Oliveira" birthdate="2010-09-23" gender="F" nation="BRA" license="403428" athleteid="1501" externalid="403428">
              <RESULTS>
                <RESULT eventid="1139" points="302" swimtime="00:01:14.86" resultid="1502" heatid="2371" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="307" swimtime="00:00:33.97" resultid="1503" heatid="2390" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Stipp Silva" birthdate="2009-12-02" gender="M" nation="BRA" license="378462" athleteid="1496" externalid="378462">
              <RESULTS>
                <RESULT eventid="1126" points="430" swimtime="00:00:59.37" resultid="1497" heatid="2369" lane="5" entrytime="00:01:00.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="336" swimtime="00:00:35.86" resultid="1498" heatid="2377" lane="4" entrytime="00:00:36.60" entrycourse="SCM" />
                <RESULT eventid="1271" points="424" swimtime="00:00:26.83" resultid="1499" heatid="2393" lane="4" entrytime="00:00:26.88" entrycourse="SCM" />
                <RESULT eventid="1457" points="344" swimtime="00:01:18.82" resultid="1500" heatid="2423" lane="5" entrytime="00:01:21.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Keirrison" lastname="Leite Silva" birthdate="2011-08-02" gender="M" nation="BRA" license="392161" athleteid="1493" externalid="392161">
              <RESULTS>
                <RESULT eventid="1178" points="100" swimtime="00:00:53.72" resultid="1494" heatid="2377" lane="7" />
                <RESULT eventid="1457" points="105" swimtime="00:01:57.13" resultid="1495" heatid="2422" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique De Oliveira" birthdate="2009-07-28" gender="M" nation="BRA" license="414505" athleteid="1488" externalid="414505">
              <RESULTS>
                <RESULT eventid="1126" points="340" swimtime="00:01:04.19" resultid="1489" heatid="2369" lane="1" entrytime="00:01:05.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1323" points="275" swimtime="00:01:13.41" resultid="1490" heatid="2401" lane="6" entrytime="00:01:14.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="341" swimtime="00:00:28.83" resultid="1491" heatid="2393" lane="7" entrytime="00:00:28.47" entrycourse="SCM" />
                <RESULT eventid="1431" points="367" swimtime="00:00:30.36" resultid="1492" heatid="2419" lane="8" entrytime="00:00:31.24" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Giroldo Santos" birthdate="2011-05-16" gender="M" nation="BRA" license="399602" athleteid="1507" externalid="399602">
              <RESULTS>
                <RESULT eventid="1323" points="126" swimtime="00:01:35.23" resultid="1508" heatid="2401" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="153" swimtime="00:00:40.58" resultid="1509" heatid="2418" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="CAMPO MOURÃO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1364" points="302" swimtime="00:04:32.26" resultid="1510" heatid="2407" lane="2" entrytime="00:04:06.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.76" />
                    <SPLIT distance="100" swimtime="00:01:00.46" />
                    <SPLIT distance="150" swimtime="00:01:35.46" />
                    <SPLIT distance="200" swimtime="00:02:15.83" />
                    <SPLIT distance="250" swimtime="00:02:49.35" />
                    <SPLIT distance="300" swimtime="00:03:27.79" />
                    <SPLIT distance="350" swimtime="00:03:57.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1496" number="1" />
                    <RELAYPOSITION athleteid="1507" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1504" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1488" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1485" points="255" swimtime="00:05:13.62" resultid="1511" heatid="2428" lane="2" entrytime="00:05:07.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.08" />
                    <SPLIT distance="100" swimtime="00:01:32.97" />
                    <SPLIT distance="150" swimtime="00:02:07.64" />
                    <SPLIT distance="200" swimtime="00:02:49.62" />
                    <SPLIT distance="250" swimtime="00:03:21.99" />
                    <SPLIT distance="300" swimtime="00:04:01.67" />
                    <SPLIT distance="350" swimtime="00:04:35.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1507" number="1" />
                    <RELAYPOSITION athleteid="1496" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1488" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1504" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="1489" nation="BRA" region="PR" clubid="1752" name="Seleção De Foz Do Iguaçu/PR" shortname="Foz Do Iguaçu">
          <ATHLETES>
            <ATHLETE firstname="Mayumi" lastname="Napole" birthdate="2010-02-01" gender="F" nation="BRA" license="376446" athleteid="1838" externalid="376446" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1284" points="307" swimtime="00:02:56.20" resultid="1839" heatid="2396" lane="8" entrytime="00:02:46.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.98" />
                    <SPLIT distance="100" swimtime="00:01:24.49" />
                    <SPLIT distance="150" swimtime="00:02:10.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="312" swimtime="00:03:18.39" resultid="1840" heatid="2387" lane="7" entrytime="00:03:17.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.26" />
                    <SPLIT distance="100" swimtime="00:01:32.58" />
                    <SPLIT distance="150" swimtime="00:02:24.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="315" swimtime="00:01:20.66" resultid="1841" heatid="2408" lane="5" entrytime="00:01:17.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1444" points="330" swimtime="00:01:30.21" resultid="1842" heatid="2420" lane="4" entrytime="00:01:28.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ysadora" lastname="Bertoldo" birthdate="2010-04-09" gender="F" nation="BRA" license="376444" athleteid="1811" externalid="376444" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1061" points="462" swimtime="00:19:34.38" resultid="1812" heatid="2359" lane="5" entrytime="00:19:50.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                    <SPLIT distance="100" swimtime="00:01:13.84" />
                    <SPLIT distance="150" swimtime="00:01:52.12" />
                    <SPLIT distance="200" swimtime="00:02:30.20" />
                    <SPLIT distance="250" swimtime="00:03:08.12" />
                    <SPLIT distance="300" swimtime="00:03:46.46" />
                    <SPLIT distance="350" swimtime="00:04:25.19" />
                    <SPLIT distance="400" swimtime="00:05:03.66" />
                    <SPLIT distance="450" swimtime="00:05:42.33" />
                    <SPLIT distance="500" swimtime="00:06:21.11" />
                    <SPLIT distance="550" swimtime="00:07:00.22" />
                    <SPLIT distance="600" swimtime="00:07:39.86" />
                    <SPLIT distance="650" swimtime="00:08:19.37" />
                    <SPLIT distance="700" swimtime="00:08:58.28" />
                    <SPLIT distance="750" swimtime="00:09:37.68" />
                    <SPLIT distance="800" swimtime="00:10:17.10" />
                    <SPLIT distance="850" swimtime="00:10:57.04" />
                    <SPLIT distance="900" swimtime="00:11:36.64" />
                    <SPLIT distance="950" swimtime="00:12:17.39" />
                    <SPLIT distance="1000" swimtime="00:12:57.47" />
                    <SPLIT distance="1050" swimtime="00:13:38.03" />
                    <SPLIT distance="1100" swimtime="00:14:17.97" />
                    <SPLIT distance="1150" swimtime="00:14:57.93" />
                    <SPLIT distance="1200" swimtime="00:15:38.08" />
                    <SPLIT distance="1250" swimtime="00:16:18.40" />
                    <SPLIT distance="1300" swimtime="00:16:58.89" />
                    <SPLIT distance="1350" swimtime="00:17:39.03" />
                    <SPLIT distance="1400" swimtime="00:18:18.66" />
                    <SPLIT distance="1450" swimtime="00:18:58.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1284" points="318" swimtime="00:02:54.14" resultid="1813" heatid="2396" lane="1" entrytime="00:02:45.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.26" />
                    <SPLIT distance="100" swimtime="00:01:26.21" />
                    <SPLIT distance="150" swimtime="00:02:11.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="436" swimtime="00:05:04.84" resultid="1814" heatid="2383" lane="2" entrytime="00:05:01.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                    <SPLIT distance="100" swimtime="00:01:14.18" />
                    <SPLIT distance="150" swimtime="00:01:52.44" />
                    <SPLIT distance="200" swimtime="00:02:31.35" />
                    <SPLIT distance="250" swimtime="00:03:10.26" />
                    <SPLIT distance="300" swimtime="00:03:48.69" />
                    <SPLIT distance="350" swimtime="00:04:27.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="442" swimtime="00:02:24.74" resultid="1815" heatid="2413" lane="6" entrytime="00:02:24.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                    <SPLIT distance="100" swimtime="00:01:10.77" />
                    <SPLIT distance="150" swimtime="00:01:48.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Marques Petry" birthdate="2008-01-08" gender="M" nation="BRA" license="392351" athleteid="1791" externalid="392351" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1152" points="276" swimtime="00:02:44.02" resultid="1792" heatid="2374" lane="8" entrytime="00:02:55.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                    <SPLIT distance="100" swimtime="00:01:16.97" />
                    <SPLIT distance="150" swimtime="00:02:01.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="426" swimtime="00:04:42.01" resultid="1793" heatid="2385" lane="1" entrytime="00:04:42.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.83" />
                    <SPLIT distance="100" swimtime="00:01:05.04" />
                    <SPLIT distance="150" swimtime="00:01:41.37" />
                    <SPLIT distance="200" swimtime="00:02:18.40" />
                    <SPLIT distance="250" swimtime="00:02:55.13" />
                    <SPLIT distance="300" swimtime="00:03:31.27" />
                    <SPLIT distance="350" swimtime="00:04:07.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="272" swimtime="00:11:19.14" resultid="1794" heatid="2425" lane="4" entrytime="00:10:13.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                    <SPLIT distance="100" swimtime="00:01:11.53" />
                    <SPLIT distance="150" swimtime="00:01:50.02" />
                    <SPLIT distance="200" swimtime="00:02:29.84" />
                    <SPLIT distance="250" swimtime="00:03:09.73" />
                    <SPLIT distance="300" swimtime="00:03:52.26" />
                    <SPLIT distance="350" swimtime="00:04:36.71" />
                    <SPLIT distance="400" swimtime="00:05:21.94" />
                    <SPLIT distance="450" swimtime="00:06:05.69" />
                    <SPLIT distance="500" swimtime="00:06:50.90" />
                    <SPLIT distance="550" swimtime="00:07:36.25" />
                    <SPLIT distance="600" swimtime="00:08:23.15" />
                    <SPLIT distance="650" swimtime="00:09:08.83" />
                    <SPLIT distance="700" swimtime="00:09:52.65" />
                    <SPLIT distance="750" swimtime="00:10:36.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1405" points="379" swimtime="00:02:17.22" resultid="1795" heatid="2415" lane="8" entrytime="00:02:19.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                    <SPLIT distance="100" swimtime="00:01:05.13" />
                    <SPLIT distance="150" swimtime="00:01:41.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Rogge" birthdate="2008-09-02" gender="M" nation="BRA" license="383387" athleteid="1763" externalid="383387" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1126" points="424" swimtime="00:00:59.66" resultid="1764" heatid="2370" lane="2" entrytime="00:00:55.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="376" swimtime="00:02:31.88" resultid="1765" heatid="2360" lane="5" entrytime="00:02:42.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                    <SPLIT distance="100" swimtime="00:01:11.81" />
                    <SPLIT distance="150" swimtime="00:01:57.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="469" swimtime="00:00:25.94" resultid="1766" heatid="2394" lane="2" entrytime="00:00:25.67" entrycourse="SCM" />
                <RESULT eventid="1431" points="381" swimtime="00:00:29.99" resultid="1767" heatid="2418" lane="2" entrytime="00:00:36.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Marques Petry" birthdate="2008-01-08" gender="M" nation="BRA" license="392352" athleteid="1796" externalid="392352" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1245" points="324" swimtime="00:02:54.90" resultid="1797" heatid="2388" lane="4" entrytime="00:03:02.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.55" />
                    <SPLIT distance="100" swimtime="00:01:24.75" />
                    <SPLIT distance="150" swimtime="00:02:10.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" status="RJC" swimtime="00:00:00.00" resultid="1798" entrytime="00:05:03.43" entrycourse="SCM" />
                <RESULT eventid="1349" points="347" swimtime="00:05:33.91" resultid="1799" heatid="2405" lane="7" entrytime="00:05:37.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                    <SPLIT distance="100" swimtime="00:01:15.30" />
                    <SPLIT distance="150" swimtime="00:02:00.17" />
                    <SPLIT distance="200" swimtime="00:02:45.01" />
                    <SPLIT distance="250" swimtime="00:03:33.49" />
                    <SPLIT distance="300" swimtime="00:04:20.99" />
                    <SPLIT distance="350" swimtime="00:04:57.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" points="332" swimtime="00:01:19.78" resultid="1800" heatid="2423" lane="6" entrytime="00:01:22.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Marques Lima" birthdate="2010-04-30" gender="F" nation="BRA" license="383051" athleteid="1824" externalid="383051">
              <RESULTS>
                <RESULT eventid="1113" points="346" swimtime="00:00:35.95" resultid="1825" heatid="2366" lane="5" entrytime="00:00:40.00" entrycourse="SCM" />
                <RESULT eventid="1284" points="348" swimtime="00:02:49.05" resultid="1826" heatid="2395" lane="3" entrytime="00:02:50.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.41" />
                    <SPLIT distance="100" swimtime="00:01:21.39" />
                    <SPLIT distance="150" swimtime="00:02:05.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="329" swimtime="00:01:19.46" resultid="1827" heatid="2408" lane="6" entrytime="00:01:18.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Faisal" lastname="Basem Ghotme" birthdate="2010-12-18" gender="M" nation="BRA" license="390809" athleteid="1843" externalid="390809" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1100" points="419" swimtime="00:00:29.54" resultid="1844" heatid="2365" lane="3" entrytime="00:00:30.57" entrycourse="SCM" />
                <RESULT eventid="1297" points="368" swimtime="00:02:27.30" resultid="1845" heatid="2398" lane="3" entrytime="00:02:25.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.35" />
                    <SPLIT distance="100" swimtime="00:01:11.72" />
                    <SPLIT distance="150" swimtime="00:01:50.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="365" swimtime="00:00:28.19" resultid="1846" heatid="2394" lane="1" entrytime="00:00:26.32" entrycourse="SCM" />
                <RESULT eventid="1379" points="396" swimtime="00:01:05.81" resultid="1847" heatid="2411" lane="8" entrytime="00:01:08.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luisa" lastname="Franco" birthdate="2010-06-09" gender="F" nation="BRA" license="383849" athleteid="1768" externalid="383849">
              <RESULTS>
                <RESULT eventid="1310" points="370" swimtime="00:01:15.28" resultid="1769" heatid="2399" lane="4" entrytime="00:01:25.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1418" points="410" swimtime="00:00:32.80" resultid="1770" heatid="2416" lane="4" entrytime="00:00:37.01" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Carvalho Carelli" birthdate="2011-10-15" gender="M" nation="BRA" license="403146" athleteid="1828" externalid="403146" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1152" points="276" swimtime="00:02:44.01" resultid="1829" heatid="2374" lane="7" entrytime="00:02:53.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                    <SPLIT distance="100" swimtime="00:01:16.75" />
                    <SPLIT distance="150" swimtime="00:02:01.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1323" points="332" swimtime="00:01:08.94" resultid="1830" heatid="2401" lane="5" entrytime="00:01:10.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1405" points="357" swimtime="00:02:19.95" resultid="1831" heatid="2415" lane="1" entrytime="00:02:19.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.26" />
                    <SPLIT distance="100" swimtime="00:01:08.06" />
                    <SPLIT distance="150" swimtime="00:01:44.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="340" swimtime="00:00:31.14" resultid="1832" heatid="2418" lane="4" entrytime="00:00:32.78" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Leticia Sbardelatti" birthdate="2011-07-28" gender="F" nation="BRA" license="403147" athleteid="1801" externalid="403147" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1139" points="284" swimtime="00:01:16.41" resultid="1802" heatid="2371" lane="7" entrytime="00:01:16.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" status="DSQ" swimtime="00:00:00.00" resultid="1803" heatid="2379" lane="2" entrytime="00:00:46.32" entrycourse="SCM" />
                <RESULT eventid="1258" points="313" swimtime="00:00:33.75" resultid="1804" heatid="2390" lane="5" entrytime="00:00:35.18" entrycourse="SCM" />
                <RESULT eventid="1418" points="213" swimtime="00:00:40.79" resultid="1805" heatid="2416" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Targat Pinheiro" birthdate="2008-09-04" gender="F" nation="BRA" license="331610" athleteid="1753" externalid="331610" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1165" points="371" swimtime="00:02:46.43" resultid="1754" heatid="2375" lane="5" entrytime="00:03:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.98" />
                    <SPLIT distance="100" swimtime="00:01:16.93" />
                    <SPLIT distance="150" swimtime="00:02:02.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="455" swimtime="00:02:38.39" resultid="1755" heatid="2363" lane="2" entrytime="00:02:43.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                    <SPLIT distance="100" swimtime="00:01:13.19" />
                    <SPLIT distance="150" swimtime="00:02:01.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="449" swimtime="00:01:10.55" resultid="1756" heatid="2400" lane="5" entrytime="00:01:12.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1418" points="476" swimtime="00:00:31.21" resultid="1757" heatid="2417" lane="3" entrytime="00:00:32.51" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Resende Ames" birthdate="2010-02-02" gender="M" nation="BRA" license="365505" athleteid="1833" externalid="365505" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1126" points="424" swimtime="00:00:59.66" resultid="1834" heatid="2369" lane="4" entrytime="00:00:59.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="427" swimtime="00:02:20.25" resultid="1835" heatid="2398" lane="4" entrytime="00:02:19.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                    <SPLIT distance="100" swimtime="00:01:07.33" />
                    <SPLIT distance="150" swimtime="00:01:43.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="397" swimtime="00:01:05.75" resultid="1836" heatid="2411" lane="3" entrytime="00:01:05.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="356" swimtime="00:00:30.67" resultid="1837" heatid="2418" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Carolina Ghellere" birthdate="2007-06-05" gender="F" nation="BRA" license="312662" athleteid="1758" externalid="312662" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1165" points="561" swimtime="00:02:25.01" resultid="1759" heatid="2376" lane="4" entrytime="00:02:26.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                    <SPLIT distance="100" swimtime="00:01:08.83" />
                    <SPLIT distance="150" swimtime="00:01:46.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="616" swimtime="00:04:31.76" resultid="1760" heatid="2383" lane="5" entrytime="00:04:51.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                    <SPLIT distance="100" swimtime="00:01:04.72" />
                    <SPLIT distance="150" swimtime="00:01:38.18" />
                    <SPLIT distance="200" swimtime="00:02:12.54" />
                    <SPLIT distance="250" swimtime="00:02:46.76" />
                    <SPLIT distance="300" swimtime="00:03:21.57" />
                    <SPLIT distance="350" swimtime="00:03:57.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1336" points="521" swimtime="00:05:21.77" resultid="1761" heatid="2403" lane="4" entrytime="00:05:25.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                    <SPLIT distance="100" swimtime="00:01:10.74" />
                    <SPLIT distance="150" swimtime="00:01:54.74" />
                    <SPLIT distance="200" swimtime="00:02:36.98" />
                    <SPLIT distance="250" swimtime="00:03:22.35" />
                    <SPLIT distance="300" swimtime="00:04:08.42" />
                    <SPLIT distance="350" swimtime="00:04:45.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="621" swimtime="00:02:09.29" resultid="1762" heatid="2413" lane="4" entrytime="00:02:11.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.29" />
                    <SPLIT distance="100" swimtime="00:01:02.09" />
                    <SPLIT distance="150" swimtime="00:01:35.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabrizzio" lastname="Paolo Cazzola" birthdate="2009-06-15" gender="M" nation="BRA" license="357168" athleteid="1786" externalid="357168" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1074" points="331" swimtime="00:02:38.42" resultid="1787" heatid="2360" lane="4" entrytime="00:02:36.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                    <SPLIT distance="100" swimtime="00:01:13.89" />
                    <SPLIT distance="150" swimtime="00:02:03.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="314" swimtime="00:02:35.34" resultid="1788" heatid="2398" lane="7" entrytime="00:02:32.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.64" />
                    <SPLIT distance="100" swimtime="00:01:16.09" />
                    <SPLIT distance="150" swimtime="00:01:56.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="374" swimtime="00:04:54.53" resultid="1789" heatid="2384" lane="6" entrytime="00:05:15.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.06" />
                    <SPLIT distance="100" swimtime="00:01:08.93" />
                    <SPLIT distance="150" swimtime="00:01:46.21" />
                    <SPLIT distance="200" swimtime="00:02:23.77" />
                    <SPLIT distance="250" swimtime="00:03:02.27" />
                    <SPLIT distance="300" swimtime="00:03:41.10" />
                    <SPLIT distance="350" swimtime="00:04:19.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1379" points="322" swimtime="00:01:10.51" resultid="1790" heatid="2410" lane="5" entrytime="00:01:09.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Geórgia" lastname="Adeli Jesus" birthdate="2008-03-27" gender="F" nation="BRA" license="312649" athleteid="1816" externalid="312649">
              <RESULTS>
                <RESULT eventid="1061" points="356" swimtime="00:21:21.38" resultid="1817" heatid="2359" lane="6" entrytime="00:21:19.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.25" />
                    <SPLIT distance="100" swimtime="00:01:14.41" />
                    <SPLIT distance="150" swimtime="00:01:54.10" />
                    <SPLIT distance="200" swimtime="00:02:35.10" />
                    <SPLIT distance="250" swimtime="00:03:16.76" />
                    <SPLIT distance="300" swimtime="00:03:58.40" />
                    <SPLIT distance="350" swimtime="00:04:40.08" />
                    <SPLIT distance="400" swimtime="00:05:22.90" />
                    <SPLIT distance="450" swimtime="00:06:06.18" />
                    <SPLIT distance="500" swimtime="00:06:49.21" />
                    <SPLIT distance="550" swimtime="00:07:32.68" />
                    <SPLIT distance="600" swimtime="00:08:15.94" />
                    <SPLIT distance="650" swimtime="00:08:59.64" />
                    <SPLIT distance="700" swimtime="00:09:43.64" />
                    <SPLIT distance="750" swimtime="00:10:27.00" />
                    <SPLIT distance="800" swimtime="00:11:10.25" />
                    <SPLIT distance="850" swimtime="00:11:53.92" />
                    <SPLIT distance="900" swimtime="00:12:38.23" />
                    <SPLIT distance="950" swimtime="00:13:22.49" />
                    <SPLIT distance="1000" swimtime="00:14:06.32" />
                    <SPLIT distance="1050" swimtime="00:14:50.70" />
                    <SPLIT distance="1100" swimtime="00:15:35.23" />
                    <SPLIT distance="1150" swimtime="00:16:19.87" />
                    <SPLIT distance="1200" swimtime="00:17:03.58" />
                    <SPLIT distance="1250" swimtime="00:17:47.83" />
                    <SPLIT distance="1300" swimtime="00:18:30.94" />
                    <SPLIT distance="1350" swimtime="00:19:14.36" />
                    <SPLIT distance="1400" swimtime="00:19:57.43" />
                    <SPLIT distance="1450" swimtime="00:20:39.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="410" swimtime="00:05:11.15" resultid="1818" heatid="2383" lane="8" entrytime="00:05:11.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.95" />
                    <SPLIT distance="100" swimtime="00:01:13.00" />
                    <SPLIT distance="150" swimtime="00:01:51.86" />
                    <SPLIT distance="200" swimtime="00:02:31.94" />
                    <SPLIT distance="250" swimtime="00:03:12.11" />
                    <SPLIT distance="300" swimtime="00:03:52.86" />
                    <SPLIT distance="350" swimtime="00:04:33.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1392" points="396" swimtime="00:02:30.14" resultid="1819" heatid="2413" lane="5" entrytime="00:02:24.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.64" />
                    <SPLIT distance="100" swimtime="00:01:10.95" />
                    <SPLIT distance="150" swimtime="00:01:49.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Christopher" lastname="De Araujo" birthdate="2008-08-09" gender="M" nation="BRA" license="366376" athleteid="1771" externalid="366376" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1245" points="422" swimtime="00:02:40.09" resultid="1772" heatid="2389" lane="2" entrytime="00:02:40.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                    <SPLIT distance="100" swimtime="00:01:16.52" />
                    <SPLIT distance="150" swimtime="00:01:58.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="489" swimtime="00:04:57.85" resultid="1773" heatid="2405" lane="2" entrytime="00:05:05.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.20" />
                    <SPLIT distance="100" swimtime="00:01:08.94" />
                    <SPLIT distance="150" swimtime="00:01:48.12" />
                    <SPLIT distance="200" swimtime="00:02:26.17" />
                    <SPLIT distance="250" swimtime="00:03:09.13" />
                    <SPLIT distance="300" swimtime="00:03:52.60" />
                    <SPLIT distance="350" swimtime="00:04:26.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="565" swimtime="00:08:52.66" resultid="1774" heatid="2426" lane="7" entrytime="00:09:14.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.43" />
                    <SPLIT distance="100" swimtime="00:01:01.68" />
                    <SPLIT distance="150" swimtime="00:01:34.72" />
                    <SPLIT distance="200" swimtime="00:02:08.05" />
                    <SPLIT distance="250" swimtime="00:02:41.43" />
                    <SPLIT distance="300" swimtime="00:03:14.93" />
                    <SPLIT distance="350" swimtime="00:03:48.75" />
                    <SPLIT distance="400" swimtime="00:04:22.62" />
                    <SPLIT distance="450" swimtime="00:04:56.21" />
                    <SPLIT distance="500" swimtime="00:05:30.29" />
                    <SPLIT distance="550" swimtime="00:06:04.68" />
                    <SPLIT distance="600" swimtime="00:06:39.03" />
                    <SPLIT distance="650" swimtime="00:07:13.05" />
                    <SPLIT distance="700" swimtime="00:07:47.49" />
                    <SPLIT distance="750" swimtime="00:08:23.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1405" points="563" swimtime="00:02:00.30" resultid="1775" heatid="2415" lane="3" entrytime="00:02:01.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.70" />
                    <SPLIT distance="100" swimtime="00:00:57.41" />
                    <SPLIT distance="150" swimtime="00:01:28.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Victoria Portela" birthdate="2009-12-04" gender="F" nation="BRA" license="383047" athleteid="1820" externalid="383047">
              <RESULTS>
                <RESULT eventid="1139" points="434" swimtime="00:01:06.33" resultid="1821" heatid="2372" lane="2" entrytime="00:01:05.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="345" swimtime="00:00:40.42" resultid="1822" heatid="2379" lane="6" entrytime="00:00:45.00" entrycourse="SCM" />
                <RESULT eventid="1258" points="468" swimtime="00:00:29.53" resultid="1823" heatid="2391" lane="4" entrytime="00:00:29.33" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Axel" lastname="Ariel Giménez González" birthdate="2011-06-01" gender="M" nation="BRA" license="365755" athleteid="1848" externalid="365755" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1126" points="394" swimtime="00:01:01.16" resultid="1849" heatid="2369" lane="2" entrytime="00:01:04.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="331" swimtime="00:00:36.05" resultid="1850" heatid="2377" lane="6" entrytime="00:00:38.67" entrycourse="SCM" />
                <RESULT eventid="1271" points="366" swimtime="00:00:28.17" resultid="1851" heatid="2393" lane="8" entrytime="00:00:29.00" entrycourse="SCM" />
                <RESULT eventid="1457" points="282" swimtime="00:01:24.22" resultid="1852" heatid="2423" lane="2" entrytime="00:01:26.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Bailke" birthdate="2007-05-04" gender="M" nation="BRA" license="370566" athleteid="1776" externalid="370566" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1152" points="230" swimtime="00:02:54.33" resultid="1777" heatid="2374" lane="1" entrytime="00:02:53.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                    <SPLIT distance="100" swimtime="00:01:17.92" />
                    <SPLIT distance="150" swimtime="00:02:04.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="300" swimtime="00:02:43.70" resultid="1778" heatid="2360" lane="3" entrytime="00:02:43.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.43" />
                    <SPLIT distance="100" swimtime="00:01:15.54" />
                    <SPLIT distance="150" swimtime="00:02:07.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1323" points="312" swimtime="00:01:10.38" resultid="1779" heatid="2401" lane="3" entrytime="00:01:11.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1470" points="344" swimtime="00:10:28.13" resultid="1780" heatid="2425" lane="5" entrytime="00:10:23.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.35" />
                    <SPLIT distance="100" swimtime="00:01:10.69" />
                    <SPLIT distance="150" swimtime="00:01:49.70" />
                    <SPLIT distance="200" swimtime="00:02:29.08" />
                    <SPLIT distance="250" swimtime="00:03:08.55" />
                    <SPLIT distance="300" swimtime="00:03:48.48" />
                    <SPLIT distance="350" swimtime="00:04:30.08" />
                    <SPLIT distance="400" swimtime="00:05:11.06" />
                    <SPLIT distance="450" swimtime="00:05:52.22" />
                    <SPLIT distance="500" swimtime="00:06:34.02" />
                    <SPLIT distance="550" swimtime="00:07:12.59" />
                    <SPLIT distance="600" swimtime="00:07:52.53" />
                    <SPLIT distance="650" swimtime="00:08:31.58" />
                    <SPLIT distance="700" swimtime="00:09:11.91" />
                    <SPLIT distance="750" swimtime="00:09:51.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanna" lastname="Mattiello" birthdate="2009-04-11" gender="F" nation="BRA" license="367011" athleteid="1781" externalid="367011" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1139" points="416" swimtime="00:01:07.31" resultid="1782" heatid="2372" lane="7" entrytime="00:01:07.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="316" swimtime="00:00:37.05" resultid="1783" heatid="2366" lane="3" entrytime="00:00:40.00" entrycourse="SCM" />
                <RESULT eventid="1258" points="411" swimtime="00:00:30.83" resultid="1784" heatid="2391" lane="6" entrytime="00:00:30.48" entrycourse="SCM" />
                <RESULT eventid="1366" points="299" swimtime="00:01:22.02" resultid="1785" heatid="2408" lane="2" entrytime="00:01:20.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Gabriel Dreher" birthdate="2011-12-05" gender="M" nation="BRA" license="403148" athleteid="1806" externalid="403148" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1100" points="202" swimtime="00:00:37.63" resultid="1807" heatid="2364" lane="5" entrytime="00:00:41.66" entrycourse="SCM" />
                <RESULT eventid="1178" points="166" swimtime="00:00:45.32" resultid="1808" heatid="2377" lane="2" entrytime="00:00:49.18" entrycourse="SCM" />
                <RESULT eventid="1323" points="126" swimtime="00:01:35.06" resultid="1809" heatid="2401" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1457" status="DSQ" swimtime="00:01:36.67" resultid="1810" heatid="2422" lane="4" entrytime="00:01:44.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="FOZ DO IGUACU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1364" points="511" swimtime="00:03:48.58" resultid="1855" heatid="2407" lane="5" entrytime="00:03:35.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.20" />
                    <SPLIT distance="100" swimtime="00:00:55.70" />
                    <SPLIT distance="150" swimtime="00:01:24.04" />
                    <SPLIT distance="200" swimtime="00:01:55.19" />
                    <SPLIT distance="250" swimtime="00:02:22.46" />
                    <SPLIT distance="300" swimtime="00:02:52.46" />
                    <SPLIT distance="350" swimtime="00:03:18.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1771" number="1" />
                    <RELAYPOSITION athleteid="1833" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1843" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1763" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1485" status="DSQ" swimtime="00:04:20.72" resultid="1856" heatid="2428" lane="5" entrytime="00:04:04.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                    <SPLIT distance="100" swimtime="00:01:05.56" />
                    <SPLIT distance="150" swimtime="00:01:39.10" />
                    <SPLIT distance="200" swimtime="00:02:18.15" />
                    <SPLIT distance="250" swimtime="00:02:48.54" />
                    <SPLIT distance="300" swimtime="00:03:24.32" />
                    <SPLIT distance="350" swimtime="00:03:50.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1843" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="1771" number="2" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION athleteid="1833" number="3" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION athleteid="1763" number="4" reactiontime="0" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="FOZ DO IGUACU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1362" points="496" swimtime="00:04:19.50" resultid="1853" heatid="2406" lane="3" entrytime="00:04:22.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                    <SPLIT distance="100" swimtime="00:01:06.37" />
                    <SPLIT distance="150" swimtime="00:01:37.75" />
                    <SPLIT distance="200" swimtime="00:02:12.39" />
                    <SPLIT distance="250" swimtime="00:02:41.57" />
                    <SPLIT distance="300" swimtime="00:03:13.21" />
                    <SPLIT distance="350" swimtime="00:03:45.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1820" number="1" />
                    <RELAYPOSITION athleteid="1753" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1758" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1811" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1483" points="435" swimtime="00:04:56.00" resultid="1854" heatid="2427" lane="5" entrytime="00:04:50.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                    <SPLIT distance="100" swimtime="00:01:18.76" />
                    <SPLIT distance="150" swimtime="00:01:56.31" />
                    <SPLIT distance="200" swimtime="00:02:40.02" />
                    <SPLIT distance="250" swimtime="00:03:11.83" />
                    <SPLIT distance="300" swimtime="00:03:51.32" />
                    <SPLIT distance="350" swimtime="00:04:21.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1811" number="1" />
                    <RELAYPOSITION athleteid="1758" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1753" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1781" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="FOZ DO IGUACU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1204" points="469" swimtime="00:02:02.41" resultid="1857" heatid="2381" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1833" number="1" />
                    <RELAYPOSITION athleteid="1771" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1758" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1753" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="1177" nation="BRA" region="PR" clubid="2048" name="Seleção De Toledo/PR" shortname="Toledo">
          <ATHLETES>
            <ATHLETE firstname="Luis" lastname="Fernando Braga Da Silva" birthdate="2011-01-10" gender="M" nation="BRA" license="380291" athleteid="2063" externalid="380291">
              <RESULTS>
                <RESULT eventid="1126" status="RJC" swimtime="00:00:00.00" resultid="2064" />
                <RESULT eventid="1100" points="213" swimtime="00:00:36.98" resultid="2065" heatid="2364" lane="3" />
                <RESULT eventid="1178" status="RJC" swimtime="00:00:00.00" resultid="2066" />
                <RESULT eventid="1271" status="RJC" swimtime="00:00:00.00" resultid="2067" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Pauly Follmann" birthdate="2011-04-19" gender="F" nation="BRA" license="413886" athleteid="2068" externalid="413886">
              <RESULTS>
                <RESULT eventid="1139" status="RJC" swimtime="00:00:00.00" resultid="2069" entrytime="00:01:34.43" entrycourse="SCM" />
                <RESULT eventid="1113" points="210" swimtime="00:00:42.44" resultid="2070" heatid="2366" lane="6" entrytime="00:00:44.59" entrycourse="SCM" />
                <RESULT eventid="1191" points="191" swimtime="00:00:49.23" resultid="2071" heatid="2379" lane="7" entrytime="00:00:50.48" entrycourse="SCM" />
                <RESULT eventid="1258" status="DSQ" swimtime="00:00:49.01" resultid="2072" heatid="2390" lane="3" entrytime="00:00:39.77" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Marafon" birthdate="2011-03-23" gender="F" nation="BRA" license="380287" swrid="5652623" athleteid="2059" externalid="380287">
              <RESULTS>
                <RESULT eventid="1191" points="399" swimtime="00:00:38.52" resultid="2060" heatid="2380" lane="6" entrytime="00:00:38.58" entrycourse="SCM" />
                <RESULT eventid="1232" points="350" swimtime="00:03:10.78" resultid="2061" heatid="2386" lane="3" entrytime="00:03:35.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.43" />
                    <SPLIT distance="100" swimtime="00:01:27.65" />
                    <SPLIT distance="150" swimtime="00:02:18.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="396" swimtime="00:00:31.22" resultid="2062" heatid="2391" lane="1" entrytime="00:00:30.93" entrycourse="SCM" />
                <RESULT eventid="1444" points="374" swimtime="00:01:26.51" resultid="2429" heatid="2421" lane="1" entrytime="00:01:24.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Welter Levandowski" birthdate="2011-05-06" gender="F" nation="BRA" license="380286" athleteid="2054" externalid="380286">
              <RESULTS>
                <RESULT eventid="1165" points="214" swimtime="00:03:19.86" resultid="2055" heatid="2375" lane="4" entrytime="00:03:13.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.49" />
                    <SPLIT distance="100" swimtime="00:01:32.82" />
                    <SPLIT distance="150" swimtime="00:02:26.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1061" points="295" swimtime="00:22:43.82" resultid="2056" heatid="2359" lane="1" entrytime="00:22:39.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:03:33.68" />
                    <SPLIT distance="100" swimtime="00:04:19.84" />
                    <SPLIT distance="150" swimtime="00:05:05.57" />
                    <SPLIT distance="200" swimtime="00:05:51.40" />
                    <SPLIT distance="250" swimtime="00:06:38.10" />
                    <SPLIT distance="300" swimtime="00:07:24.54" />
                    <SPLIT distance="350" swimtime="00:08:10.06" />
                    <SPLIT distance="400" swimtime="00:08:53.63" />
                    <SPLIT distance="450" swimtime="00:09:39.27" />
                    <SPLIT distance="500" swimtime="00:10:25.79" />
                    <SPLIT distance="550" swimtime="00:11:11.33" />
                    <SPLIT distance="600" swimtime="00:11:56.71" />
                    <SPLIT distance="650" swimtime="00:12:43.66" />
                    <SPLIT distance="700" swimtime="00:13:31.03" />
                    <SPLIT distance="750" swimtime="00:14:17.98" />
                    <SPLIT distance="800" swimtime="00:15:04.71" />
                    <SPLIT distance="850" swimtime="00:15:51.75" />
                    <SPLIT distance="900" swimtime="00:16:38.92" />
                    <SPLIT distance="950" swimtime="00:17:25.84" />
                    <SPLIT distance="1000" swimtime="00:18:12.52" />
                    <SPLIT distance="1050" swimtime="00:18:59.25" />
                    <SPLIT distance="1100" swimtime="00:19:45.21" />
                    <SPLIT distance="1150" swimtime="00:20:31.04" />
                    <SPLIT distance="1200" swimtime="00:21:15.96" />
                    <SPLIT distance="1250" swimtime="00:22:00.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="228" swimtime="00:01:28.46" resultid="2057" heatid="2399" lane="5" entrytime="00:01:26.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1206" points="340" swimtime="00:05:31.08" resultid="2058" heatid="2382" lane="3" entrytime="00:05:26.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                    <SPLIT distance="100" swimtime="00:01:16.64" />
                    <SPLIT distance="150" swimtime="00:01:57.95" />
                    <SPLIT distance="200" swimtime="00:02:40.87" />
                    <SPLIT distance="250" swimtime="00:03:23.88" />
                    <SPLIT distance="300" swimtime="00:04:07.61" />
                    <SPLIT distance="350" swimtime="00:04:50.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Torres Romancini" birthdate="2010-05-28" gender="F" nation="BRA" license="347218" athleteid="2049" externalid="347218">
              <RESULTS>
                <RESULT eventid="1113" points="439" swimtime="00:00:33.20" resultid="2050" heatid="2367" lane="6" entrytime="00:00:33.68" entrycourse="SCM" />
                <RESULT eventid="1284" points="419" swimtime="00:02:38.89" resultid="2051" heatid="2395" lane="5" entrytime="00:02:48.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.09" />
                    <SPLIT distance="100" swimtime="00:01:16.30" />
                    <SPLIT distance="150" swimtime="00:01:57.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="420" swimtime="00:01:13.25" resultid="2052" heatid="2409" lane="6" entrytime="00:01:13.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1418" points="346" swimtime="00:00:34.71" resultid="2053" heatid="2417" lane="7" entrytime="00:00:33.64" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Marafon Duarte" birthdate="2011-08-18" gender="M" nation="BRA" license="414184" athleteid="2078" externalid="414184">
              <RESULTS>
                <RESULT eventid="1126" points="213" swimtime="00:01:15.01" resultid="2079" heatid="2368" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" status="RJC" swimtime="00:00:00.00" resultid="2080" />
                <RESULT eventid="1271" points="237" swimtime="00:00:32.55" resultid="2081" heatid="2392" lane="5" />
                <RESULT eventid="1431" points="145" swimtime="00:00:41.39" resultid="2082" heatid="2418" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kawan" lastname="Gustavo Klein Ladeia" birthdate="2010-04-19" gender="M" nation="BRA" license="413943" athleteid="2073" externalid="413943">
              <RESULTS>
                <RESULT eventid="1126" status="RJC" swimtime="00:00:00.00" resultid="2074" />
                <RESULT eventid="1178" points="212" swimtime="00:00:41.78" resultid="2075" heatid="2377" lane="1" />
                <RESULT eventid="1271" status="RJC" swimtime="00:00:00.00" resultid="2076" />
                <RESULT eventid="1457" points="205" swimtime="00:01:33.61" resultid="2077" heatid="2422" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="TOLEDO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1362" points="307" swimtime="00:05:04.35" resultid="2083" heatid="2406" lane="2" entrytime="00:05:33.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="100" swimtime="00:01:07.92" />
                    <SPLIT distance="150" swimtime="00:01:39.96" />
                    <SPLIT distance="200" swimtime="00:02:17.21" />
                    <SPLIT distance="250" swimtime="00:02:51.98" />
                    <SPLIT distance="300" swimtime="00:03:31.09" />
                    <SPLIT distance="350" swimtime="00:04:19.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2059" number="1" />
                    <RELAYPOSITION athleteid="2049" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2054" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="2068" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1483" status="DSQ" swimtime="00:05:35.68" resultid="2084" heatid="2427" lane="6" entrytime="00:06:10.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                    <SPLIT distance="100" swimtime="00:01:16.47" />
                    <SPLIT distance="150" swimtime="00:01:56.12" />
                    <SPLIT distance="200" swimtime="00:02:41.43" />
                    <SPLIT distance="250" swimtime="00:03:20.58" />
                    <SPLIT distance="300" swimtime="00:04:10.96" />
                    <SPLIT distance="350" swimtime="00:04:53.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="2" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION number="3" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION number="4" reactiontime="0" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="TOLEDO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1204" points="312" swimtime="00:02:20.26" resultid="2085" heatid="2381" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                    <SPLIT distance="100" swimtime="00:01:15.68" />
                    <SPLIT distance="150" swimtime="00:01:48.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2063" number="1" />
                    <RELAYPOSITION athleteid="2059" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2049" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="2073" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="6462" nation="BRA" region="PR" clubid="2042" name="Seleção De São José Dos Pinhais/PR" shortname="São José Dos Pinhais">
          <ATHLETES>
            <ATHLETE firstname="Diego" lastname="Brasil Caropreso" birthdate="2009-10-29" gender="M" nation="BRA" license="399502" athleteid="2043" externalid="399502">
              <RESULTS>
                <RESULT eventid="1126" points="384" swimtime="00:01:01.69" resultid="2044" heatid="2369" lane="3" entrytime="00:01:03.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="304" swimtime="00:02:42.91" resultid="2045" heatid="2360" lane="2" entrytime="00:02:54.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.97" />
                    <SPLIT distance="100" swimtime="00:01:18.48" />
                    <SPLIT distance="150" swimtime="00:02:07.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1271" points="385" swimtime="00:00:27.70" resultid="2046" heatid="2393" lane="6" entrytime="00:00:28.33" entrycourse="SCM" />
                <RESULT eventid="1405" points="400" swimtime="00:02:14.77" resultid="2047" heatid="2414" lane="7" entrytime="00:02:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                    <SPLIT distance="100" swimtime="00:01:03.90" />
                    <SPLIT distance="150" swimtime="00:01:39.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
