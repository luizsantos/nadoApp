<?xml version="1.0" encoding="UTF-8"?>
<LENEX revisiondate="2024-12-02" created="2025-03-23T22:59:17" version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.81460">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Foz do Iguaçu" name="Torneio Regional da 2ª Região (Pré-Mirim/Sênior)" course="SCM" deadline="2025-03-09" entrystartdate="2025-01-27" entrytype="INVITATION" hostclub="Universidade Estadual de Maringá" hostclub.url="http://www.uem.br/" number="39515" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/evento/natacao/39515" startmethod="1" status="OFFICIAL" timing="AUTOMATIC" touchpad="ONESIDE" masters="F" withdrawuntil="2025-03-10" state="PR" nation="BRA" hytek.courseorder="S">
      <AGEDATE value="2025-03-08" type="YEAR" />
      <POOL name="Ginásio de Esportes Costa Cavalcante" lanemin="1" lanemax="6" />
      <FACILITY city="Foz do Iguaçu" name="Ginásio de Esportes Costa Cavalcante" nation="BRA" state="PR" street="Rua Lisboa, 510" street2="Jardim Alice" zip="85858-050" />
      <POINTTABLE pointtableid="3017" name="AQUA Point Scoring" version="2024" />
      <QUALIFY from="2024-03-08" until="2025-03-07" />
      <CONTACT city="Curitiba" email="ti@swimtimebrasil.com" fax="+55 (41) 99252-0598" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99252-0598" street="Avenida do Batel, 1230" street2="Sala 202" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2025-03-15" daytime="08:40" endtime="22:19" number="1" officialmeeting="08:00" status="OFFICIAL" teamleadermeeting="08:30" warmupfrom="07:30" warmupuntil="08:30">
          <EVENTS>
            <EVENT eventid="1060" daytime="08:40" gender="F" number="1" order="1" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1061" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2912" />
                    <RANKING order="2" place="2" resultid="2690" />
                    <RANKING order="3" place="3" resultid="2686" />
                    <RANKING order="4" place="4" resultid="3095" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2818" />
                    <RANKING order="2" place="2" resultid="2662" />
                    <RANKING order="3" place="3" resultid="2920" />
                    <RANKING order="4" place="4" resultid="2924" />
                    <RANKING order="5" place="5" resultid="2916" />
                    <RANKING order="6" place="6" resultid="2448" />
                    <RANKING order="7" place="7" resultid="2610" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3101" daytime="08:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3102" daytime="08:44" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1063" daytime="08:50" gender="M" number="2" order="2" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1064" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2949" />
                    <RANKING order="2" place="2" resultid="2953" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2635" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3103" daytime="08:50" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1066" daytime="08:56" gender="F" number="3" order="3" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1067" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2858" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2555" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2434" />
                    <RANKING order="2" place="2" resultid="2439" />
                    <RANKING order="3" place="3" resultid="2552" />
                    <RANKING order="4" place="4" resultid="2868" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1071" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3013" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1073" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3104" daytime="08:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3105" daytime="09:00" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1074" daytime="09:04" gender="M" number="4" order="4" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1075" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2587" />
                    <RANKING order="2" place="2" resultid="2879" />
                    <RANKING order="3" place="3" resultid="2601" />
                    <RANKING order="4" place="-1" resultid="2854" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1076" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1077" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2829" />
                    <RANKING order="2" place="2" resultid="3048" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1078" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2465" />
                    <RANKING order="2" place="2" resultid="2519" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1079" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2526" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1080" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1081" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3106" daytime="09:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3107" daytime="09:08" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1082" daytime="09:12" gender="F" number="5" order="5" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1083" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3098" />
                    <RANKING order="2" place="2" resultid="2616" />
                    <RANKING order="3" place="3" resultid="3096" />
                    <RANKING order="4" place="-1" resultid="2458" />
                    <RANKING order="5" place="-1" resultid="3036" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1084" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2947" />
                    <RANKING order="2" place="2" resultid="2450" />
                    <RANKING order="3" place="3" resultid="3092" />
                    <RANKING order="4" place="4" resultid="2584" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3108" daytime="09:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3109" daytime="09:14" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1085" daytime="09:16" gender="M" number="6" order="6" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1086" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2620" />
                    <RANKING order="2" place="2" resultid="2951" />
                    <RANKING order="3" place="3" resultid="2736" />
                    <RANKING order="4" place="4" resultid="2955" />
                    <RANKING order="5" place="5" resultid="2652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1087" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2636" />
                    <RANKING order="2" place="2" resultid="2593" />
                    <RANKING order="3" place="-1" resultid="2672" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3110" daytime="09:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3111" daytime="09:18" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1088" daytime="09:22" gender="F" number="7" order="7" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1089" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2898" />
                    <RANKING order="2" place="2" resultid="2606" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1090" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1091" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1092" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1093" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1094" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3012" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1095" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2715" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3112" daytime="09:22" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1096" daytime="09:24" gender="M" number="8" order="8" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1097" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2496" />
                    <RANKING order="2" place="2" resultid="3059" />
                    <RANKING order="3" place="3" resultid="3067" />
                    <RANKING order="4" place="-1" resultid="3063" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2540" />
                    <RANKING order="2" place="2" resultid="2490" />
                    <RANKING order="3" place="3" resultid="2999" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1099" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3047" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1100" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2464" />
                    <RANKING order="2" place="2" resultid="3021" />
                    <RANKING order="3" place="3" resultid="2482" />
                    <RANKING order="4" place="4" resultid="2536" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1101" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2514" />
                    <RANKING order="2" place="2" resultid="2479" />
                    <RANKING order="3" place="3" resultid="2722" />
                    <RANKING order="4" place="4" resultid="2874" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1103" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2461" />
                    <RANKING order="2" place="2" resultid="3008" />
                    <RANKING order="3" place="3" resultid="3026" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3113" daytime="09:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3114" daytime="09:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3115" daytime="09:28" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3116" daytime="09:30" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1104" daytime="09:32" gender="F" number="9" order="9" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1105" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2692" />
                    <RANKING order="2" place="2" resultid="3099" />
                    <RANKING order="3" place="3" resultid="3035" />
                    <RANKING order="4" place="4" resultid="3071" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1106" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2820" />
                    <RANKING order="2" place="2" resultid="2922" />
                    <RANKING order="3" place="3" resultid="2918" />
                    <RANKING order="4" place="4" resultid="2570" />
                    <RANKING order="5" place="5" resultid="2851" />
                    <RANKING order="6" place="6" resultid="2583" />
                    <RANKING order="7" place="7" resultid="2905" />
                    <RANKING order="8" place="8" resultid="3087" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3117" daytime="09:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3118" daytime="09:34" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1107" daytime="09:36" gender="M" number="10" order="10" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1108" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2619" />
                    <RANKING order="2" place="2" resultid="2667" />
                    <RANKING order="3" place="3" resultid="2684" />
                    <RANKING order="4" place="4" resultid="2735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1109" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2645" />
                    <RANKING order="2" place="2" resultid="2592" />
                    <RANKING order="3" place="3" resultid="2640" />
                    <RANKING order="4" place="4" resultid="3078" />
                    <RANKING order="5" place="5" resultid="3081" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3119" daytime="09:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3120" daytime="09:38" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1110" daytime="09:42" gender="F" number="11" order="11" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1111" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2578" />
                    <RANKING order="2" place="2" resultid="3030" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1112" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2560" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1113" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2433" />
                    <RANKING order="2" place="2" resultid="2547" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1114" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1115" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2523" />
                    <RANKING order="2" place="2" resultid="2746" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1116" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2834" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1117" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3121" daytime="09:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3122" daytime="09:44" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1118" daytime="09:48" gender="M" number="12" order="12" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1119" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2595" />
                    <RANKING order="2" place="2" resultid="3039" />
                    <RANKING order="3" place="3" resultid="2573" />
                    <RANKING order="4" place="4" resultid="2600" />
                    <RANKING order="5" place="5" resultid="2994" />
                    <RANKING order="6" place="6" resultid="3062" />
                    <RANKING order="7" place="-1" resultid="2631" />
                    <RANKING order="8" place="-1" resultid="2853" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1120" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2883" />
                    <RANKING order="2" place="2" resultid="2893" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1121" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1122" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2863" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1123" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1124" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3017" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1125" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3123" daytime="09:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3124" daytime="09:50" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1126" daytime="10:08" gender="F" number="13" order="14" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1127" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2691" />
                    <RANKING order="2" place="2" resultid="2688" />
                    <RANKING order="3" place="3" resultid="2615" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2926" />
                    <RANKING order="2" place="2" resultid="2917" />
                    <RANKING order="3" place="3" resultid="2904" />
                    <RANKING order="4" place="4" resultid="2569" />
                    <RANKING order="5" place="5" resultid="3093" />
                    <RANKING order="6" place="6" resultid="2850" />
                    <RANKING order="7" place="7" resultid="2612" />
                    <RANKING order="8" place="-1" resultid="2582" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3125" daytime="10:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3126" daytime="10:10" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1129" daytime="10:12" gender="M" number="14" order="15" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1130" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2683" />
                    <RANKING order="2" place="2" resultid="2651" />
                    <RANKING order="3" place="3" resultid="2734" />
                    <RANKING order="4" place="-1" resultid="2623" />
                    <RANKING order="5" place="-1" resultid="2954" />
                    <RANKING order="6" place="-1" resultid="2968" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1131" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2644" />
                    <RANKING order="2" place="-1" resultid="2671" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3127" daytime="10:12" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1132" daytime="10:14" gender="F" number="15" order="16" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1133" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1134" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2559" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1135" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2551" />
                    <RANKING order="2" place="2" resultid="3043" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1136" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1137" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1138" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2824" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1139" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3128" daytime="10:14" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1140" daytime="10:18" gender="M" number="16" order="17" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1141" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3058" />
                    <RANKING order="2" place="2" resultid="3061" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1142" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2474" />
                    <RANKING order="2" place="2" resultid="3053" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1143" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2453" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1144" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2518" />
                    <RANKING order="2" place="2" resultid="3003" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1145" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1146" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1147" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3007" />
                    <RANKING order="2" place="2" resultid="2564" />
                    <RANKING order="3" place="3" resultid="2648" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3129" daytime="10:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3130" daytime="10:18" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1148" daytime="10:22" gender="F" number="17" order="18" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1149" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2914" />
                    <RANKING order="2" place="2" resultid="2687" />
                    <RANKING order="3" place="3" resultid="2614" />
                    <RANKING order="4" place="4" resultid="2457" />
                    <RANKING order="5" place="5" resultid="3070" />
                    <RANKING order="6" place="6" resultid="3097" />
                    <RANKING order="7" place="7" resultid="3034" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2664" />
                    <RANKING order="2" place="2" resultid="2946" />
                    <RANKING order="3" place="3" resultid="2925" />
                    <RANKING order="4" place="4" resultid="2849" />
                    <RANKING order="5" place="5" resultid="3094" />
                    <RANKING order="6" place="6" resultid="2903" />
                    <RANKING order="7" place="7" resultid="2611" />
                    <RANKING order="8" place="8" resultid="3086" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3131" daytime="10:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3132" daytime="10:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3133" daytime="10:24" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1151" daytime="10:28" gender="M" number="18" order="19" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1152" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2618" />
                    <RANKING order="2" place="2" resultid="2666" />
                    <RANKING order="3" place="3" resultid="2950" />
                    <RANKING order="4" place="4" resultid="2682" />
                    <RANKING order="5" place="5" resultid="2622" />
                    <RANKING order="6" place="6" resultid="2650" />
                    <RANKING order="7" place="-1" resultid="2967" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1153" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2643" />
                    <RANKING order="2" place="2" resultid="2639" />
                    <RANKING order="3" place="3" resultid="2591" />
                    <RANKING order="4" place="4" resultid="3080" />
                    <RANKING order="5" place="5" resultid="3077" />
                    <RANKING order="6" place="-1" resultid="2670" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3134" daytime="10:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3135" daytime="10:28" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1154" daytime="10:32" gender="F" number="19" order="20" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1155" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2845" />
                    <RANKING order="2" place="2" resultid="2605" />
                    <RANKING order="3" place="3" resultid="3029" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1156" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2554" />
                    <RANKING order="2" place="2" resultid="2932" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1157" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2438" />
                    <RANKING order="2" place="2" resultid="2550" />
                    <RANKING order="3" place="3" resultid="3042" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1158" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2505" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1159" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2509" />
                    <RANKING order="2" place="2" resultid="2522" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1160" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2823" />
                    <RANKING order="2" place="2" resultid="3011" />
                    <RANKING order="3" place="3" resultid="2726" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1161" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2714" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3136" daytime="10:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3137" daytime="10:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3138" daytime="10:34" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1162" daytime="10:36" gender="M" number="20" order="21" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1163" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2586" />
                    <RANKING order="2" place="2" resultid="2907" />
                    <RANKING order="3" place="3" resultid="2572" />
                    <RANKING order="4" place="4" resultid="3038" />
                    <RANKING order="5" place="5" resultid="2878" />
                    <RANKING order="6" place="6" resultid="2630" />
                    <RANKING order="7" place="7" resultid="2495" />
                    <RANKING order="8" place="8" resultid="3057" />
                    <RANKING order="9" place="9" resultid="2993" />
                    <RANKING order="10" place="10" resultid="3066" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1164" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2473" />
                    <RANKING order="2" place="2" resultid="2539" />
                    <RANKING order="3" place="3" resultid="2839" />
                    <RANKING order="4" place="4" resultid="3052" />
                    <RANKING order="5" place="5" resultid="2998" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1165" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2531" />
                    <RANKING order="2" place="2" resultid="2452" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1166" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3020" />
                    <RANKING order="2" place="2" resultid="3002" />
                    <RANKING order="3" place="3" resultid="2535" />
                    <RANKING order="4" place="4" resultid="3073" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1167" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2478" />
                    <RANKING order="2" place="2" resultid="2721" />
                    <RANKING order="3" place="3" resultid="2873" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1168" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2428" />
                    <RANKING order="2" place="2" resultid="3016" />
                    <RANKING order="3" place="3" resultid="2717" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1169" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3006" />
                    <RANKING order="2" place="2" resultid="3025" />
                    <RANKING order="3" place="3" resultid="2647" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3139" daytime="10:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3140" daytime="10:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3141" daytime="10:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3142" daytime="10:42" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3143" daytime="10:44" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1170" daytime="10:46" gender="F" number="21" order="22" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1171" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3465" />
                    <RANKING order="2" place="2" resultid="3464" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1172" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3419" />
                    <RANKING order="2" place="2" resultid="3353" />
                    <RANKING order="3" place="3" resultid="3495" />
                    <RANKING order="4" place="4" resultid="3447" />
                    <RANKING order="5" place="5" resultid="3247" />
                    <RANKING order="6" place="6" resultid="3366" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1173" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3430" />
                    <RANKING order="2" place="2" resultid="3286" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1174" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1175" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3323" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1176" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1177" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1178" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1179" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3144" daytime="10:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3145" daytime="10:50" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1180" daytime="10:54" gender="M" number="22" order="23" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1181" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3313" />
                    <RANKING order="2" place="2" resultid="3374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1182" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3378" />
                    <RANKING order="2" place="2" resultid="3277" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1183" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3297" />
                    <RANKING order="2" place="2" resultid="3506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1184" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3483" />
                    <RANKING order="2" place="2" resultid="3244" />
                    <RANKING order="3" place="-1" resultid="3399" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1185" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3336" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1187" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3348" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1188" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3258" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1189" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3402" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3146" daytime="10:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3147" daytime="11:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3148" daytime="11:04" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1190" daytime="11:08" gender="F" number="23" order="24" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1191" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3499" />
                    <RANKING order="2" place="2" resultid="3448" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1192" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3436" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1193" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3452" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1194" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1195" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1196" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3471" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1197" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3149" daytime="11:08" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1198" daytime="11:34" gender="M" number="24" order="25" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1199" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1200" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3468" />
                    <RANKING order="2" place="2" resultid="3496" />
                    <RANKING order="3" place="3" resultid="3502" />
                    <RANKING order="4" place="-1" resultid="3484" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1201" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3433" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1202" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3439" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1203" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3262" />
                    <RANKING order="2" place="2" resultid="3301" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1204" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1205" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3150" daytime="11:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3151" daytime="12:00" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2025-03-15" daytime="15:40" endtime="13:22" number="2" officialmeeting="15:00" status="OFFICIAL" teamleadermeeting="15:30" warmupfrom="14:30" warmupuntil="15:30">
          <EVENTS>
            <EVENT eventid="1206" daytime="15:40" gender="F" number="25" order="1" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1207" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="1208" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3310" />
                    <RANKING order="2" place="2" resultid="3427" />
                    <RANKING order="3" place="3" resultid="3389" />
                    <RANKING order="4" place="4" resultid="3359" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3152" daytime="15:40" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1209" daytime="15:44" gender="M" number="26" order="2" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1210" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3317" />
                    <RANKING order="2" place="2" resultid="3488" />
                    <RANKING order="3" place="3" resultid="3474" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1211" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3407" />
                    <RANKING order="2" place="2" resultid="3477" />
                    <RANKING order="3" place="3" resultid="3424" />
                    <RANKING order="4" place="4" resultid="3414" />
                    <RANKING order="5" place="-1" resultid="3252" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3153" daytime="15:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3154" daytime="15:46" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1212" daytime="15:50" gender="F" number="27" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1213" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1214" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1215" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1216" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1217" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1218" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1219" agemax="-1" agemin="20" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1220" daytime="15:50" gender="M" number="28" order="4" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1221" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3456" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1222" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3485" />
                    <RANKING order="2" place="-1" resultid="3503" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1223" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3338" />
                    <RANKING order="2" place="2" resultid="3434" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1224" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1225" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3263" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1226" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1227" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3155" daytime="15:50" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1228" daytime="15:58" gender="F" number="29" order="5" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1229" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3370" />
                    <RANKING order="2" place="2" resultid="3344" />
                    <RANKING order="3" place="3" resultid="3332" />
                    <RANKING order="4" place="4" resultid="3306" />
                    <RANKING order="5" place="5" resultid="3292" />
                    <RANKING order="6" place="6" resultid="3272" />
                    <RANKING order="7" place="7" resultid="3329" />
                    <RANKING order="8" place="8" resultid="3357" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3156" daytime="15:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3157" daytime="15:58" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1230" daytime="16:00" gender="M" number="30" order="6" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1231" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3375" />
                    <RANKING order="2" place="2" resultid="3320" />
                    <RANKING order="3" place="3" resultid="3266" />
                    <RANKING order="4" place="4" resultid="3396" />
                    <RANKING order="5" place="5" resultid="3340" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3158" daytime="16:00" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1232" daytime="16:02" gender="F" number="31" order="7" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1233" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3480" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1234" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3428" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3159" daytime="16:02" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1235" daytime="16:06" gender="M" number="32" order="8" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1236" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3318" />
                    <RANKING order="2" place="2" resultid="3255" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1237" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3283" />
                    <RANKING order="2" place="2" resultid="3478" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3160" daytime="16:06" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1238" daytime="16:08" gender="F" number="33" order="9" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1239" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1240" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3438" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1241" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3250" />
                    <RANKING order="2" place="2" resultid="3248" />
                    <RANKING order="3" place="-1" resultid="3453" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1242" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1243" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3410" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1244" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3472" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1245" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3161" daytime="16:08" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1246" daytime="16:16" gender="M" number="34" order="10" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1247" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3299" />
                    <RANKING order="2" place="2" resultid="3382" />
                    <RANKING order="3" place="3" resultid="3422" />
                    <RANKING order="4" place="-1" resultid="3463" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1248" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3470" />
                    <RANKING order="2" place="2" resultid="3498" />
                    <RANKING order="3" place="3" resultid="3245" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1249" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3365" />
                    <RANKING order="2" place="2" resultid="3513" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1250" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3405" />
                    <RANKING order="2" place="2" resultid="3441" />
                    <RANKING order="3" place="3" resultid="3372" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1251" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1252" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1253" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3162" daytime="16:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3163" daytime="16:24" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1254" daytime="16:32" gender="F" number="35" order="11" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1255" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3442" />
                    <RANKING order="2" place="2" resultid="3314" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1256" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3311" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3164" daytime="16:32" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1257" daytime="16:34" gender="M" number="36" order="12" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1258" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="1259" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3425" />
                    <RANKING order="2" place="2" resultid="3408" />
                    <RANKING order="3" place="3" resultid="3392" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3165" daytime="16:34" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1260" daytime="16:36" gender="F" number="37" order="13" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1261" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1262" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1263" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1264" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1265" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1266" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3420" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1267" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3166" daytime="16:36" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1268" daytime="16:40" gender="M" number="38" order="14" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1269" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3347" />
                    <RANKING order="2" place="2" resultid="3380" />
                    <RANKING order="3" place="3" resultid="3423" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1270" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3504" />
                    <RANKING order="2" place="-1" resultid="3486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1271" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3241" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1272" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3406" />
                    <RANKING order="2" place="2" resultid="3373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1273" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3350" />
                    <RANKING order="2" place="2" resultid="3445" />
                    <RANKING order="3" place="-1" resultid="3379" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1274" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3260" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1275" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3167" daytime="16:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3168" daytime="16:42" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1276" daytime="16:46" gender="F" number="39" order="15" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1277" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3369" />
                    <RANKING order="2" place="2" resultid="3331" />
                    <RANKING order="3" place="3" resultid="3343" />
                    <RANKING order="4" place="4" resultid="3291" />
                    <RANKING order="5" place="5" resultid="3305" />
                    <RANKING order="6" place="6" resultid="3328" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3169" daytime="16:46" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1278" daytime="16:48" gender="M" number="40" order="16" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1279" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3376" />
                    <RANKING order="2" place="2" resultid="3397" />
                    <RANKING order="3" place="3" resultid="3267" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3170" daytime="16:48" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1280" daytime="17:04" gender="F" number="41" order="18" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1281" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3270" />
                    <RANKING order="2" place="2" resultid="3315" />
                    <RANKING order="3" place="3" resultid="3443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1282" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3390" />
                    <RANKING order="2" place="2" resultid="3295" />
                    <RANKING order="3" place="3" resultid="3360" />
                    <RANKING order="4" place="4" resultid="3387" />
                    <RANKING order="5" place="5" resultid="3281" />
                    <RANKING order="6" place="6" resultid="3510" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3171" daytime="17:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3172" daytime="17:06" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1283" daytime="17:08" gender="M" number="42" order="19" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1284" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3319" />
                    <RANKING order="2" place="2" resultid="3256" />
                    <RANKING order="3" place="3" resultid="3475" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1285" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3479" />
                    <RANKING order="2" place="2" resultid="3274" />
                    <RANKING order="3" place="3" resultid="3393" />
                    <RANKING order="4" place="4" resultid="3354" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3173" daytime="17:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3174" daytime="17:12" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1286" daytime="17:14" gender="F" number="43" order="20" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1287" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3287" />
                    <RANKING order="2" place="2" resultid="3524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1288" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3362" />
                    <RANKING order="2" place="-1" resultid="3412" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1289" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3324" />
                    <RANKING order="2" place="2" resultid="3528" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1290" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1291" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3278" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1292" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3473" />
                    <RANKING order="2" place="2" resultid="3308" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1293" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3175" daytime="17:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3176" daytime="17:16" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1294" daytime="17:18" gender="M" number="44" order="21" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1295" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3327" />
                    <RANKING order="2" place="2" resultid="3521" />
                    <RANKING order="3" place="-1" resultid="3383" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1296" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3304" />
                    <RANKING order="2" place="2" resultid="3517" />
                    <RANKING order="3" place="3" resultid="3526" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1297" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1298" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3523" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1299" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1300" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3508" />
                    <RANKING order="2" place="2" resultid="3418" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1301" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3403" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3177" daytime="17:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3178" daytime="17:22" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1302" daytime="17:24" gender="F" number="45" order="22" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1303" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3307" />
                    <RANKING order="2" place="2" resultid="3273" />
                    <RANKING order="3" place="3" resultid="3330" />
                    <RANKING order="4" place="4" resultid="3358" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3179" daytime="17:24" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1304" daytime="17:26" gender="M" number="46" order="23" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1305" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3341" />
                    <RANKING order="2" place="2" resultid="3321" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3180" daytime="17:26" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1306" daytime="17:28" gender="F" number="47" order="24" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1307" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3269" />
                    <RANKING order="2" place="2" resultid="3459" />
                    <RANKING order="3" place="3" resultid="3493" />
                    <RANKING order="4" place="4" resultid="3457" />
                    <RANKING order="5" place="5" resultid="3481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1308" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3312" />
                    <RANKING order="2" place="2" resultid="3294" />
                    <RANKING order="3" place="3" resultid="3429" />
                    <RANKING order="4" place="4" resultid="3386" />
                    <RANKING order="5" place="5" resultid="3491" />
                    <RANKING order="6" place="6" resultid="3280" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3181" daytime="17:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3182" daytime="17:30" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1309" daytime="17:34" gender="M" number="48" order="25" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1310" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3257" />
                    <RANKING order="2" place="2" resultid="3489" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1311" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3284" />
                    <RANKING order="2" place="2" resultid="3415" />
                    <RANKING order="3" place="3" resultid="3275" />
                    <RANKING order="4" place="4" resultid="3466" />
                    <RANKING order="5" place="5" resultid="3355" />
                    <RANKING order="6" place="-1" resultid="3253" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3183" daytime="17:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3184" daytime="17:36" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1312" daytime="17:38" gender="F" number="49" order="26" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1313" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3431" />
                    <RANKING order="2" place="2" resultid="3501" />
                    <RANKING order="3" place="3" resultid="3449" />
                    <RANKING order="4" place="4" resultid="3351" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1314" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1315" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1316" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1317" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1318" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3505" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1319" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3185" daytime="17:38" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1320" daytime="17:42" gender="M" number="50" order="27" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1321" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3290" />
                    <RANKING order="2" place="-1" resultid="3381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1322" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3401" />
                    <RANKING order="2" place="2" resultid="3246" />
                    <RANKING order="3" place="-1" resultid="3335" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1323" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3435" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1324" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3515" />
                    <RANKING order="2" place="2" resultid="3368" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1325" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3302" />
                    <RANKING order="2" place="2" resultid="3264" />
                    <RANKING order="3" place="3" resultid="3446" />
                    <RANKING order="4" place="4" resultid="3385" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1326" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3243" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1327" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3300" />
                    <RANKING order="2" place="2" resultid="3507" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3186" daytime="17:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3187" daytime="17:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3188" daytime="17:46" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1328" daytime="17:50" gender="F" number="51" order="28" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1329" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3371" />
                    <RANKING order="2" place="2" resultid="3345" />
                    <RANKING order="3" place="3" resultid="3333" />
                    <RANKING order="4" place="4" resultid="3293" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3189" daytime="17:50" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1330" daytime="17:52" gender="M" number="52" order="29" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1331" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3398" />
                    <RANKING order="2" place="2" resultid="3377" />
                    <RANKING order="3" place="3" resultid="3268" />
                    <RANKING order="4" place="4" resultid="3322" />
                    <RANKING order="5" place="5" resultid="3342" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3190" daytime="17:52" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1332" daytime="17:54" gender="F" number="53" order="30" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1333" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3271" />
                    <RANKING order="2" place="2" resultid="3316" />
                    <RANKING order="3" place="3" resultid="3460" />
                    <RANKING order="4" place="4" resultid="3494" />
                    <RANKING order="5" place="5" resultid="3444" />
                    <RANKING order="6" place="6" resultid="3458" />
                    <RANKING order="7" place="7" resultid="3482" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1334" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3391" />
                    <RANKING order="2" place="2" resultid="3492" />
                    <RANKING order="3" place="3" resultid="3388" />
                    <RANKING order="4" place="4" resultid="3511" />
                    <RANKING order="5" place="5" resultid="3296" />
                    <RANKING order="6" place="6" resultid="3361" />
                    <RANKING order="7" place="7" resultid="3282" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3191" daytime="17:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3192" daytime="17:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3193" daytime="17:58" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1335" daytime="18:00" gender="M" number="54" order="31" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1336" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3490" />
                    <RANKING order="2" place="2" resultid="3476" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1337" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3285" />
                    <RANKING order="2" place="2" resultid="3409" />
                    <RANKING order="3" place="3" resultid="3276" />
                    <RANKING order="4" place="4" resultid="3416" />
                    <RANKING order="5" place="5" resultid="3426" />
                    <RANKING order="6" place="6" resultid="3467" />
                    <RANKING order="7" place="7" resultid="3394" />
                    <RANKING order="8" place="8" resultid="3356" />
                    <RANKING order="9" place="-1" resultid="3254" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3194" daytime="18:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3195" daytime="18:02" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1338" daytime="18:06" gender="F" number="55" order="32" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1339" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3432" />
                    <RANKING order="2" place="2" resultid="3288" />
                    <RANKING order="3" place="3" resultid="3352" />
                    <RANKING order="4" place="4" resultid="3525" />
                    <RANKING order="5" place="-1" resultid="3450" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1340" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3363" />
                    <RANKING order="2" place="-1" resultid="3413" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1341" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3249" />
                    <RANKING order="2" place="2" resultid="3251" />
                    <RANKING order="3" place="3" resultid="3529" />
                    <RANKING order="4" place="-1" resultid="3454" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1342" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3404" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1343" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3411" />
                    <RANKING order="2" place="2" resultid="3339" />
                    <RANKING order="3" place="3" resultid="3279" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1344" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3421" />
                    <RANKING order="2" place="2" resultid="3309" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1345" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3196" daytime="18:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3197" daytime="18:08" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3198" daytime="18:10" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1346" daytime="18:12" gender="M" number="56" order="33" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1347" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3346" />
                    <RANKING order="2" place="2" resultid="3298" />
                    <RANKING order="3" place="3" resultid="3326" />
                    <RANKING order="4" place="4" resultid="3289" />
                    <RANKING order="5" place="5" resultid="3520" />
                    <RANKING order="6" place="6" resultid="3527" />
                    <RANKING order="7" place="7" resultid="3509" />
                    <RANKING order="8" place="-1" resultid="3455" />
                    <RANKING order="9" place="-1" resultid="3462" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1348" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3303" />
                    <RANKING order="2" place="2" resultid="3469" />
                    <RANKING order="3" place="3" resultid="3497" />
                    <RANKING order="4" place="4" resultid="3400" />
                    <RANKING order="5" place="5" resultid="3516" />
                    <RANKING order="6" place="-1" resultid="3334" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1349" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3337" />
                    <RANKING order="2" place="2" resultid="3364" />
                    <RANKING order="3" place="3" resultid="3240" />
                    <RANKING order="4" place="4" resultid="3512" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1350" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3514" />
                    <RANKING order="2" place="2" resultid="3440" />
                    <RANKING order="3" place="3" resultid="3518" />
                    <RANKING order="4" place="4" resultid="3522" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1351" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3395" />
                    <RANKING order="2" place="2" resultid="3384" />
                    <RANKING order="3" place="3" resultid="3349" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1352" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3242" />
                    <RANKING order="2" place="2" resultid="3259" />
                    <RANKING order="3" place="3" resultid="3417" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1353" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3519" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3199" daytime="18:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3200" daytime="18:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3201" daytime="18:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3202" daytime="18:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3203" daytime="18:22" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3225" daytime="18:24" gender="M" number="101" order="34" round="TIMETRIAL" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3233" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3261" />
                    <RANKING order="2" place="-1" resultid="3487" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3530" daytime="18:24" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3234" daytime="18:28" gender="F" number="102" order="35" round="TIMETRIAL" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3235" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3325" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3754" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3236" daytime="18:28" gender="M" number="103" order="36" round="TIMETRIAL" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3237" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3265" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3531" daytime="18:28" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3238" daytime="18:32" gender="F" number="104" order="37" round="TIMETRIAL" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3239" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3451" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3532" daytime="18:32" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="1035" nation="BRA" region="PR" clubid="2991" swrid="93778" name="Fundação De Esportes De Campo Mourão" shortname="Fecam">
          <ATHLETES>
            <ATHLETE firstname="Fabricio" lastname="Campos Faria" birthdate="2013-09-15" gender="M" nation="BRA" license="422156" athleteid="3079" externalid="422156">
              <RESULTS>
                <RESULT eventid="1151" points="146" swimtime="00:00:38.28" resultid="3080" heatid="3134" lane="5" />
                <RESULT eventid="1107" points="68" reactiontime="+72" swimtime="00:00:54.04" resultid="3081" heatid="3119" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Ferreira Batista" birthdate="2014-11-26" gender="F" nation="BRA" license="392160" swrid="5515815" athleteid="3033" externalid="392160">
              <RESULTS>
                <RESULT eventid="1148" points="122" swimtime="00:00:46.13" resultid="3034" heatid="3132" lane="1" entrytime="00:00:42.40" entrycourse="SCM" />
                <RESULT eventid="1104" points="117" swimtime="00:00:51.61" resultid="3035" heatid="3118" lane="1" entrytime="00:00:41.83" entrycourse="SCM" />
                <RESULT comment="SW 7.1 - Mais de uma pernada de borboleta antes da primeira pernada de peito após o início ou a virada.  (Horário: 9:23), Após a volta dos 25m." eventid="1082" status="DSQ" swimtime="00:00:58.36" resultid="3036" heatid="3108" lane="4" entrytime="00:00:58.93" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Gomes De Souza" birthdate="2006-01-30" gender="F" nation="BRA" license="308464" swrid="5603844" athleteid="3010" externalid="308464">
              <RESULTS>
                <RESULT eventid="1154" points="301" swimtime="00:00:34.20" resultid="3011" heatid="3137" lane="5" entrytime="00:00:33.70" entrycourse="SCM" />
                <RESULT eventid="1088" points="242" swimtime="00:00:45.52" resultid="3012" heatid="3112" lane="2" entrytime="00:00:43.19" entrycourse="SCM" />
                <RESULT eventid="1066" points="227" swimtime="00:03:00.65" resultid="3013" heatid="3104" lane="4" entrytime="00:02:49.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                    <SPLIT distance="100" swimtime="00:01:20.87" />
                    <SPLIT distance="150" swimtime="00:02:10.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="224" swimtime="00:01:42.61" resultid="3505" heatid="3185" lane="5" entrytime="00:01:39.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rebecca" lastname="Rosasantos" birthdate="2013-01-21" gender="F" nation="BRA" license="422158" athleteid="3085" externalid="422158">
              <RESULTS>
                <RESULT eventid="1148" points="86" swimtime="00:00:51.76" resultid="3086" heatid="3131" lane="2" />
                <RESULT eventid="1104" points="58" swimtime="00:01:05.04" resultid="3087" heatid="3117" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Samuel" lastname="Massuda Santos" birthdate="2012-06-09" gender="M" nation="BRA" license="392189" swrid="5603872" athleteid="3037" externalid="392189">
              <RESULTS>
                <RESULT eventid="1162" points="250" swimtime="00:00:32.00" resultid="3038" heatid="3140" lane="4" entrytime="00:00:33.01" entrycourse="SCM" />
                <RESULT eventid="1118" points="246" reactiontime="+73" swimtime="00:01:17.09" resultid="3039" heatid="3123" lane="3" entrytime="00:01:23.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="227" swimtime="00:02:59.61" resultid="3506" heatid="3146" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaue" lastname="Guilherme Chagas" birthdate="2005-06-29" gender="M" nation="BRA" license="378464" swrid="5603851" athleteid="3024" externalid="378464">
              <RESULTS>
                <RESULT eventid="1162" points="330" swimtime="00:00:29.16" resultid="3025" heatid="3142" lane="4" entrytime="00:00:28.54" entrycourse="SCM" />
                <RESULT eventid="1096" points="243" swimtime="00:00:39.93" resultid="3026" heatid="3115" lane="6" entrytime="00:00:38.78" entrycourse="SCM" />
                <RESULT eventid="1320" points="225" swimtime="00:01:30.85" resultid="3507" heatid="3187" lane="6" entrytime="00:01:26.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Batinga Ponchielli" birthdate="2007-01-18" gender="M" nation="BRA" license="378461" swrid="5251143" athleteid="3015" externalid="378461">
              <RESULTS>
                <RESULT eventid="1162" points="318" swimtime="00:00:29.52" resultid="3016" heatid="3142" lane="2" entrytime="00:00:28.90" entrycourse="SCM" />
                <RESULT eventid="1118" points="276" swimtime="00:01:14.22" resultid="3017" heatid="3124" lane="6" entrytime="00:01:15.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1294" points="242" reactiontime="+70" swimtime="00:00:35.45" resultid="3508" heatid="3178" lane="2" entrytime="00:00:35.13" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anthony" lastname="Lira Gordo" birthdate="2012-04-09" gender="M" nation="BRA" license="415261" swrid="5757893" athleteid="3065" externalid="415261">
              <RESULTS>
                <RESULT eventid="1162" points="121" swimtime="00:00:40.65" resultid="3066" heatid="3139" lane="6" />
                <RESULT eventid="1096" points="108" swimtime="00:00:52.28" resultid="3067" heatid="3113" lane="2" />
                <RESULT eventid="1346" points="117" swimtime="00:01:31.48" resultid="3509" heatid="3199" lane="2" entrytime="00:01:34.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonia" lastname="Giglini Zambon" birthdate="2015-05-25" gender="F" nation="BRA" license="422157" athleteid="3082" externalid="422157">
              <RESULTS>
                <RESULT eventid="1280" points="40" reactiontime="+74" swimtime="00:01:13.44" resultid="3510" heatid="3172" lane="1" />
                <RESULT eventid="1332" points="87" swimtime="00:00:51.66" resultid="3511" heatid="3192" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stela" lastname="Gouveia" birthdate="2014-02-27" gender="F" nation="BRA" license="415498" swrid="5757891" athleteid="3069" externalid="415498">
              <RESULTS>
                <RESULT eventid="1148" points="130" swimtime="00:00:45.22" resultid="3070" heatid="3131" lane="3" entrytime="00:00:51.45" entrycourse="SCM" />
                <RESULT eventid="1104" points="116" reactiontime="+89" swimtime="00:00:51.66" resultid="3071" heatid="3117" lane="1" entrytime="00:00:55.31" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kenzo" lastname="Kimura" birthdate="2010-04-23" gender="M" nation="BRA" license="403429" swrid="5676289" athleteid="3046" externalid="403429">
              <RESULTS>
                <RESULT eventid="1096" points="198" swimtime="00:00:42.76" resultid="3047" heatid="3114" lane="2" entrytime="00:00:42.06" entrycourse="SCM" />
                <RESULT eventid="1074" points="226" swimtime="00:02:43.08" resultid="3048" heatid="3107" lane="1" entrytime="00:02:45.20" entrycourse="SCM" />
                <RESULT eventid="1346" points="264" swimtime="00:01:09.81" resultid="3512" heatid="3200" lane="2" entrytime="00:01:12.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1246" points="197" swimtime="00:06:04.33" resultid="3513" heatid="3162" lane="2" entrytime="00:06:26.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:16.09" />
                    <SPLIT distance="150" swimtime="00:02:00.30" />
                    <SPLIT distance="350" swimtime="00:05:14.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Stipp Silva" birthdate="2009-12-02" gender="M" nation="BRA" license="378462" swrid="5603918" athleteid="3019" externalid="378462">
              <RESULTS>
                <RESULT eventid="1162" points="469" swimtime="00:00:25.94" resultid="3020" heatid="3143" lane="1" entrytime="00:00:26.12" entrycourse="SCM" />
                <RESULT eventid="1096" points="407" swimtime="00:00:33.66" resultid="3021" heatid="3115" lane="4" entrytime="00:00:34.47" entrycourse="SCM" />
                <RESULT eventid="1346" points="463" swimtime="00:00:57.92" resultid="3514" heatid="3202" lane="3" entrytime="00:00:59.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="409" swimtime="00:01:14.44" resultid="3515" heatid="3187" lane="4" entrytime="00:01:17.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Eduardo Schork Filho" birthdate="2012-12-28" gender="M" nation="BRA" license="413906" swrid="5755352" athleteid="3056" externalid="413906">
              <RESULTS>
                <RESULT eventid="1162" points="149" swimtime="00:00:38.01" resultid="3057" heatid="3139" lane="3" entrytime="00:00:40.03" entrycourse="SCM" />
                <RESULT eventid="1140" points="128" swimtime="00:00:43.05" resultid="3058" heatid="3129" lane="2" entrytime="00:00:45.84" entrycourse="SCM" />
                <RESULT eventid="1096" points="126" swimtime="00:00:49.71" resultid="3059" heatid="3114" lane="1" entrytime="00:00:49.71" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur" lastname="Setsuo Iechika" birthdate="2013-03-10" gender="M" nation="BRA" license="422155" athleteid="3076" externalid="422155">
              <RESULTS>
                <RESULT eventid="1151" points="85" swimtime="00:00:45.74" resultid="3077" heatid="3134" lane="1" />
                <RESULT eventid="1107" points="75" reactiontime="+102" swimtime="00:00:52.39" resultid="3078" heatid="3119" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Giroldo Santos" birthdate="2011-05-16" gender="M" nation="BRA" license="399602" swrid="5755354" athleteid="3051" externalid="399602">
              <RESULTS>
                <RESULT eventid="1162" points="191" swimtime="00:00:34.95" resultid="3052" heatid="3140" lane="1" entrytime="00:00:34.40" entrycourse="SCM" />
                <RESULT eventid="1140" points="160" reactiontime="+852" swimtime="00:00:40.03" resultid="3053" heatid="3129" lane="4" entrytime="00:00:40.47" entrycourse="SCM" />
                <RESULT eventid="1346" points="195" swimtime="00:01:17.28" resultid="3516" heatid="3200" lane="5" entrytime="00:01:17.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1294" points="130" reactiontime="+82" swimtime="00:00:43.63" resultid="3517" heatid="3178" lane="1" entrytime="00:00:43.79" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique De Oliveira" birthdate="2009-07-28" gender="M" nation="BRA" license="414505" swrid="5755355" athleteid="3001" externalid="414505">
              <RESULTS>
                <RESULT eventid="1162" points="369" swimtime="00:00:28.10" resultid="3002" heatid="3143" lane="6" entrytime="00:00:27.76" entrycourse="SCM" />
                <RESULT eventid="1140" points="392" swimtime="00:00:29.71" resultid="3003" heatid="3130" lane="5" entrytime="00:00:30.11" entrycourse="SCM" />
                <RESULT eventid="1346" points="361" swimtime="00:01:02.96" resultid="3518" heatid="3202" lane="1" entrytime="00:01:04.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Franco Santos" birthdate="2002-01-03" gender="M" nation="BRA" license="290441" swrid="5546064" athleteid="3005" externalid="290441">
              <RESULTS>
                <RESULT eventid="1162" points="535" swimtime="00:00:24.83" resultid="3006" heatid="3143" lane="3" entrytime="00:00:25.20" entrycourse="SCM" />
                <RESULT eventid="1140" points="499" swimtime="00:00:27.42" resultid="3007" heatid="3130" lane="3" entrytime="00:00:27.37" entrycourse="SCM" />
                <RESULT eventid="1096" points="457" swimtime="00:00:32.39" resultid="3008" heatid="3116" lane="5" entrytime="00:00:32.25" entrycourse="SCM" />
                <RESULT eventid="1346" points="449" swimtime="00:00:58.54" resultid="3519" heatid="3203" lane="5" entrytime="00:00:56.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Franca Rebollo" birthdate="2012-09-26" gender="M" nation="BRA" license="385780" swrid="5538081" athleteid="2992" externalid="385780">
              <RESULTS>
                <RESULT eventid="1162" points="146" swimtime="00:00:38.24" resultid="2993" heatid="3139" lane="2" entrytime="00:00:40.78" entrycourse="SCM" />
                <RESULT eventid="1118" points="124" swimtime="00:01:36.77" resultid="2994" heatid="3123" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1346" points="145" swimtime="00:01:25.17" resultid="3520" heatid="3199" lane="3" entrytime="00:01:29.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1294" points="123" reactiontime="+83" swimtime="00:00:44.39" resultid="3521" heatid="3177" lane="3" entrytime="00:00:47.68" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Capel Adelino" birthdate="2009-04-24" gender="M" nation="BRA" license="422154" athleteid="3072" externalid="422154">
              <RESULTS>
                <RESULT eventid="1162" points="226" swimtime="00:00:33.06" resultid="3073" heatid="3139" lane="1" />
                <RESULT eventid="1346" points="163" swimtime="00:01:21.93" resultid="3522" heatid="3199" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1294" points="117" reactiontime="+114" swimtime="00:00:45.11" resultid="3523" heatid="3177" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Ferreira Batista" birthdate="2012-03-29" gender="F" nation="BRA" license="385779" swrid="5532525" athleteid="3028" externalid="385779">
              <RESULTS>
                <RESULT eventid="1154" points="277" swimtime="00:00:35.16" resultid="3029" heatid="3137" lane="1" entrytime="00:00:34.46" entrycourse="SCM" />
                <RESULT eventid="1110" points="239" reactiontime="+78" swimtime="00:01:28.35" resultid="3030" heatid="3121" lane="4" entrytime="00:01:33.62" entrycourse="SCM" />
                <RESULT eventid="1286" points="255" reactiontime="+63" swimtime="00:00:39.77" resultid="3524" heatid="3175" lane="3" entrytime="00:00:40.97" />
                <RESULT eventid="1338" points="258" swimtime="00:01:18.89" resultid="3525" heatid="3197" lane="6" entrytime="00:01:18.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Keirrison" lastname="Leite Silva" birthdate="2011-08-02" gender="M" nation="BRA" license="392161" swrid="5603864" athleteid="2997" externalid="392161">
              <RESULTS>
                <RESULT eventid="1162" points="150" swimtime="00:00:37.90" resultid="2998" heatid="3139" lane="4" entrytime="00:00:40.07" entrycourse="SCM" />
                <RESULT eventid="1096" points="135" swimtime="00:00:48.60" resultid="2999" heatid="3113" lane="3" entrytime="00:00:53.72" entrycourse="SCM" />
                <RESULT eventid="1294" points="81" reactiontime="+92" swimtime="00:00:50.91" resultid="3526" heatid="3177" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henry" lastname="Sadao Da Silva" birthdate="2012-10-02" gender="M" nation="BRA" license="413907" swrid="5755359" athleteid="3060" externalid="413907">
              <RESULTS>
                <RESULT eventid="1140" points="71" swimtime="00:00:52.30" resultid="3061" heatid="3129" lane="5" entrytime="00:00:52.88" entrycourse="SCM" />
                <RESULT eventid="1118" points="80" reactiontime="+74" swimtime="00:01:51.97" resultid="3062" heatid="3123" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.57" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 9:32), Na volta dos 25m." eventid="1096" status="DSQ" swimtime="00:00:55.47" resultid="3063" heatid="3113" lane="4" entrytime="00:00:59.07" entrycourse="SCM" />
                <RESULT eventid="1346" points="118" swimtime="00:01:31.26" resultid="3527" heatid="3199" lane="5" entrytime="00:01:39.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Gabrieli Oliveira" birthdate="2010-09-23" gender="F" nation="BRA" license="403428" swrid="5676288" athleteid="3041" externalid="403428">
              <RESULTS>
                <RESULT eventid="1154" points="293" swimtime="00:00:34.49" resultid="3042" heatid="3137" lane="4" entrytime="00:00:33.32" entrycourse="SCM" />
                <RESULT eventid="1132" points="238" swimtime="00:00:39.31" resultid="3043" heatid="3128" lane="1" entrytime="00:00:39.82" entrycourse="SCM" />
                <RESULT eventid="1286" points="220" reactiontime="+86" swimtime="00:00:41.78" resultid="3528" heatid="3176" lane="1" entrytime="00:00:40.96" />
                <RESULT eventid="1338" points="265" swimtime="00:01:18.23" resultid="3529" heatid="3197" lane="5" entrytime="00:01:14.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2416" nation="BRA" region="PR" clubid="2459" swrid="93758" name="Apan/Maringá">
          <ATHLETES>
            <ATHLETE firstname="Matheus" lastname="Junio Brambilla" birthdate="2002-04-08" gender="M" nation="BRA" license="392112" swrid="5603859" athleteid="2646" externalid="392112">
              <RESULTS>
                <RESULT eventid="1162" points="239" swimtime="00:00:32.46" resultid="2647" heatid="3140" lane="3" entrytime="00:00:31.73" entrycourse="SCM" />
                <RESULT eventid="1140" points="289" swimtime="00:00:32.86" resultid="2648" heatid="3130" lane="6" entrytime="00:00:31.80" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Forti Francisco" birthdate="2015-07-08" gender="M" nation="BRA" license="392104" swrid="5534395" athleteid="2625" externalid="392104">
              <RESULTS>
                <RESULT eventid="1209" status="DNS" swimtime="00:00:00.00" resultid="3252" heatid="3154" lane="3" late="yes" entrytime="00:01:33.39" />
                <RESULT eventid="1309" status="DNS" swimtime="00:00:00.00" resultid="3253" heatid="3184" lane="4" late="yes" entrytime="00:00:56.39" />
                <RESULT eventid="1335" status="DNS" swimtime="00:00:00.00" resultid="3254" heatid="3195" lane="2" late="yes" entrytime="00:00:41.32" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laion" lastname="Miguel Simoes" birthdate="2016-04-02" gender="M" nation="BRA" license="407179" swrid="5718695" athleteid="2701" externalid="407179">
              <RESULTS>
                <RESULT eventid="1235" points="93" swimtime="00:01:48.47" resultid="3255" heatid="3160" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1283" points="71" reactiontime="+78" swimtime="00:00:53.36" resultid="3256" heatid="3174" lane="5" entrytime="00:00:53.32" />
                <RESULT eventid="1309" points="84" swimtime="00:00:56.85" resultid="3257" heatid="3184" lane="1" entrytime="00:01:02.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Pacheco" birthdate="2006-12-20" gender="M" nation="BRA" license="336850" swrid="5603854" athleteid="2499" externalid="336850">
              <RESULTS>
                <RESULT eventid="1074" points="482" swimtime="00:02:06.67" resultid="2500" heatid="3107" lane="4" entrytime="00:02:09.31" entrycourse="SCM" />
                <RESULT eventid="1180" points="439" swimtime="00:02:24.23" resultid="3258" heatid="3146" lane="4" />
                <RESULT eventid="1346" points="451" swimtime="00:00:58.45" resultid="3259" heatid="3203" lane="6" entrytime="00:00:59.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="383" swimtime="00:01:05.79" resultid="3260" heatid="3168" lane="4" entrytime="00:01:02.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3225" points="428" swimtime="00:02:21.76" resultid="3261" heatid="3530" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                    <SPLIT distance="100" swimtime="00:01:08.22" />
                    <SPLIT distance="150" swimtime="00:01:45.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Da Cateburcio" birthdate="2004-01-18" gender="F" nation="BRA" license="407186" swrid="5737919" athleteid="2713" externalid="407186">
              <RESULTS>
                <RESULT eventid="1154" points="83" swimtime="00:00:52.45" resultid="2714" heatid="3136" lane="3" entrytime="00:00:52.12" entrycourse="SCM" />
                <RESULT eventid="1088" points="35" swimtime="00:01:26.27" resultid="2715" heatid="3112" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Garcia Cavalcante" birthdate="2008-08-11" gender="M" nation="BRA" license="369676" swrid="5603841" athleteid="2485" externalid="369676">
              <RESULTS>
                <RESULT eventid="1198" points="377" swimtime="00:19:31.67" resultid="3262" heatid="3151" lane="3" entrytime="00:19:37.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                    <SPLIT distance="100" swimtime="00:01:13.97" />
                    <SPLIT distance="150" swimtime="00:01:53.31" />
                    <SPLIT distance="200" swimtime="00:02:32.18" />
                    <SPLIT distance="250" swimtime="00:03:09.76" />
                    <SPLIT distance="300" swimtime="00:03:47.94" />
                    <SPLIT distance="350" swimtime="00:04:27.23" />
                    <SPLIT distance="400" swimtime="00:05:06.49" />
                    <SPLIT distance="450" swimtime="00:05:45.91" />
                    <SPLIT distance="500" swimtime="00:06:24.90" />
                    <SPLIT distance="550" swimtime="00:07:04.09" />
                    <SPLIT distance="600" swimtime="00:07:43.74" />
                    <SPLIT distance="650" swimtime="00:08:22.84" />
                    <SPLIT distance="700" swimtime="00:09:01.55" />
                    <SPLIT distance="750" swimtime="00:09:41.04" />
                    <SPLIT distance="800" swimtime="00:10:19.70" />
                    <SPLIT distance="850" swimtime="00:10:58.23" />
                    <SPLIT distance="900" swimtime="00:11:36.90" />
                    <SPLIT distance="950" swimtime="00:12:15.51" />
                    <SPLIT distance="1000" swimtime="00:12:54.43" />
                    <SPLIT distance="1050" swimtime="00:13:33.43" />
                    <SPLIT distance="1100" swimtime="00:14:12.48" />
                    <SPLIT distance="1150" swimtime="00:14:52.15" />
                    <SPLIT distance="1200" swimtime="00:15:31.77" />
                    <SPLIT distance="1250" swimtime="00:16:11.49" />
                    <SPLIT distance="1300" swimtime="00:16:51.71" />
                    <SPLIT distance="1350" swimtime="00:17:32.38" />
                    <SPLIT distance="1400" swimtime="00:18:13.14" />
                    <SPLIT distance="1450" swimtime="00:18:52.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" points="344" swimtime="00:05:34.97" resultid="3263" heatid="3155" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.69" />
                    <SPLIT distance="100" swimtime="00:01:21.85" />
                    <SPLIT distance="150" swimtime="00:02:06.05" />
                    <SPLIT distance="200" swimtime="00:02:51.13" />
                    <SPLIT distance="250" swimtime="00:03:34.95" />
                    <SPLIT distance="300" swimtime="00:04:19.20" />
                    <SPLIT distance="350" swimtime="00:04:58.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="362" swimtime="00:01:17.55" resultid="3264" heatid="3188" lane="6" entrytime="00:01:13.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3236" points="359" swimtime="00:02:48.92" resultid="3265" heatid="3531" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                    <SPLIT distance="100" swimtime="00:01:22.08" />
                    <SPLIT distance="150" swimtime="00:02:04.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Tomazeli" birthdate="2017-11-30" gender="M" nation="BRA" license="421901" athleteid="2750" externalid="421901">
              <RESULTS>
                <RESULT eventid="1230" points="26" swimtime="00:00:33.04" resultid="3266" heatid="3158" lane="4" />
                <RESULT eventid="1278" points="34" swimtime="00:00:31.54" resultid="3267" heatid="3170" lane="3" />
                <RESULT eventid="1330" points="40" swimtime="00:00:58.84" resultid="3268" heatid="3190" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Siqueira Almeida" birthdate="2016-06-21" gender="F" nation="BRA" license="414848" swrid="5755360" athleteid="2729" externalid="414848">
              <RESULTS>
                <RESULT eventid="1306" points="90" swimtime="00:01:03.15" resultid="3269" heatid="3182" lane="2" entrytime="00:01:07.24" />
                <RESULT eventid="1280" points="133" reactiontime="+63" swimtime="00:00:49.40" resultid="3270" heatid="3172" lane="3" entrytime="00:00:52.59" />
                <RESULT eventid="1332" points="106" swimtime="00:00:48.34" resultid="3271" heatid="3193" lane="3" entrytime="00:00:56.36" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luara" lastname="Polizeli Marostica" birthdate="2017-04-12" gender="F" nation="BRA" license="421958" athleteid="2805" externalid="421958">
              <RESULTS>
                <RESULT eventid="1228" points="28" swimtime="00:00:36.60" resultid="3272" heatid="3156" lane="2" />
                <RESULT eventid="1302" points="45" swimtime="00:00:36.95" resultid="3273" heatid="3179" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heitor" lastname="Bello Paula" birthdate="2015-06-14" gender="M" nation="BRA" license="393776" swrid="5507529" athleteid="2657" externalid="393776">
              <RESULTS>
                <RESULT eventid="1283" points="98" reactiontime="+67" swimtime="00:00:47.86" resultid="3274" heatid="3174" lane="4" entrytime="00:00:46.58" />
                <RESULT eventid="1309" points="89" swimtime="00:00:55.85" resultid="3275" heatid="3184" lane="5" entrytime="00:00:56.87" />
                <RESULT eventid="1335" points="134" swimtime="00:00:39.35" resultid="3276" heatid="3195" lane="4" entrytime="00:00:40.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Vaneti Mazuti" birthdate="2014-11-29" gender="M" nation="BRA" license="414850" swrid="5757897" athleteid="2733" externalid="414850">
              <RESULTS>
                <RESULT eventid="1129" points="70" swimtime="00:00:52.71" resultid="2734" heatid="3127" lane="1" entrytime="00:00:55.94" entrycourse="SCM" />
                <RESULT eventid="1107" points="92" reactiontime="+65" swimtime="00:00:48.85" resultid="2735" heatid="3119" lane="3" />
                <RESULT eventid="1085" points="109" swimtime="00:00:52.15" resultid="2736" heatid="3110" lane="3" entrytime="00:00:51.55" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Tomazeli" birthdate="2013-02-05" gender="M" nation="BRA" license="392109" swrid="5614097" athleteid="2638" externalid="392109">
              <RESULTS>
                <RESULT eventid="1151" points="226" swimtime="00:00:33.07" resultid="2639" heatid="3135" lane="2" entrytime="00:00:34.94" entrycourse="SCM" />
                <RESULT eventid="1107" points="164" reactiontime="+78" swimtime="00:00:40.37" resultid="2640" heatid="3120" lane="1" entrytime="00:00:43.14" entrycourse="SCM" />
                <RESULT eventid="1180" points="185" swimtime="00:03:12.14" resultid="3277" heatid="3147" lane="5" entrytime="00:03:22.01" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Lopes Ferreira" birthdate="2008-12-03" gender="F" nation="ESP" license="383455" athleteid="2745" externalid="383455">
              <RESULTS>
                <RESULT eventid="1110" points="254" reactiontime="+74" swimtime="00:01:26.58" resultid="2746" heatid="3121" lane="2" entrytime="00:01:35.28" entrycourse="SCM" />
                <RESULT eventid="1066" points="303" swimtime="00:02:44.13" resultid="2747" heatid="3104" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                    <SPLIT distance="150" swimtime="00:02:00.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="261" reactiontime="+75" swimtime="00:00:39.48" resultid="3278" heatid="3175" lane="2" />
                <RESULT eventid="1338" points="291" swimtime="00:01:15.80" resultid="3279" heatid="3196" lane="2" entrytime="00:01:21.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Coleto Arcanjo" birthdate="2015-08-17" gender="F" nation="BRA" license="407176" swrid="5631404" athleteid="2693" externalid="407176">
              <RESULTS>
                <RESULT eventid="1306" points="31" swimtime="00:01:29.64" resultid="3280" heatid="3182" lane="6" entrytime="00:01:18.10" />
                <RESULT eventid="1280" points="60" reactiontime="+68" swimtime="00:01:04.30" resultid="3281" heatid="3172" lane="2" entrytime="00:01:07.52" />
                <RESULT eventid="1332" points="57" swimtime="00:00:59.33" resultid="3282" heatid="3193" lane="1" entrytime="00:01:04.15" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Arthur Da Silva Ortiz" birthdate="2015-04-20" gender="M" nation="BRA" license="399733" swrid="5676285" athleteid="2673" externalid="399733">
              <RESULTS>
                <RESULT eventid="1235" points="141" swimtime="00:01:34.56" resultid="3283" heatid="3160" lane="4" entrytime="00:01:53.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1309" points="117" swimtime="00:00:50.96" resultid="3284" heatid="3184" lane="3" entrytime="00:00:48.59" />
                <RESULT eventid="1335" points="145" swimtime="00:00:38.31" resultid="3285" heatid="3195" lane="3" entrytime="00:00:39.01" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Pavão" birthdate="2012-04-04" gender="F" nation="BRA" license="377259" swrid="5603888" athleteid="2576" externalid="377259">
              <RESULTS>
                <RESULT eventid="1110" points="296" reactiontime="+59" swimtime="00:01:22.36" resultid="2578" heatid="3122" lane="5" entrytime="00:01:22.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="308" swimtime="00:03:00.25" resultid="3286" heatid="3145" lane="6" entrytime="00:03:19.45" />
                <RESULT eventid="1286" points="305" reactiontime="+61" swimtime="00:00:37.50" resultid="3287" heatid="3176" lane="2" entrytime="00:00:38.37" />
                <RESULT eventid="1338" points="314" swimtime="00:01:13.91" resultid="3288" heatid="3196" lane="4" entrytime="00:01:19.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Diogo" lastname="Sanchez" birthdate="2012-11-29" gender="M" nation="BRA" license="370658" swrid="5603906" athleteid="2494" externalid="370658">
              <RESULTS>
                <RESULT eventid="1162" points="152" swimtime="00:00:37.76" resultid="2495" heatid="3140" lane="6" entrytime="00:00:36.70" entrycourse="SCM" />
                <RESULT eventid="1096" points="206" swimtime="00:00:42.24" resultid="2496" heatid="3114" lane="5" entrytime="00:00:44.88" entrycourse="SCM" />
                <RESULT eventid="1346" points="177" swimtime="00:01:19.77" resultid="3289" heatid="3200" lane="6" entrytime="00:01:27.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="214" swimtime="00:01:32.38" resultid="3290" heatid="3186" lane="2" entrytime="00:01:39.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Fernanda Silva Simoes" birthdate="2017-09-05" gender="F" nation="BRA" license="421904" athleteid="2762" externalid="421904">
              <RESULTS>
                <RESULT eventid="1276" points="58" swimtime="00:00:30.56" resultid="3291" heatid="3169" lane="4" />
                <RESULT eventid="1228" points="32" swimtime="00:00:35.15" resultid="3292" heatid="3157" lane="3" />
                <RESULT eventid="1328" points="36" swimtime="00:01:09.33" resultid="3293" heatid="3189" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="De Araujo" birthdate="2015-08-09" gender="F" nation="BRA" license="407185" swrid="5725999" athleteid="2709" externalid="407185">
              <RESULTS>
                <RESULT eventid="1306" points="118" swimtime="00:00:57.79" resultid="3294" heatid="3182" lane="5" entrytime="00:01:07.36" />
                <RESULT eventid="1280" points="78" reactiontime="+94" swimtime="00:00:59.09" resultid="3295" heatid="3172" lane="4" entrytime="00:01:01.07" />
                <RESULT eventid="1332" points="85" reactiontime="+218" swimtime="00:00:52.01" resultid="3296" heatid="3193" lane="4" entrytime="00:00:57.05" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Ayres" birthdate="2012-05-05" gender="M" nation="BRA" license="378035" swrid="5208079" athleteid="2594" externalid="378035">
              <RESULTS>
                <RESULT eventid="1118" points="301" reactiontime="+77" swimtime="00:01:12.08" resultid="2595" heatid="3124" lane="2" entrytime="00:01:14.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="300" swimtime="00:02:43.75" resultid="3297" heatid="3148" lane="5" entrytime="00:02:49.52" />
                <RESULT eventid="1346" points="311" swimtime="00:01:06.12" resultid="3298" heatid="3201" lane="2" entrytime="00:01:05.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1246" points="353" swimtime="00:05:00.32" resultid="3299" heatid="3163" lane="5" entrytime="00:05:16.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                    <SPLIT distance="100" swimtime="00:01:10.54" />
                    <SPLIT distance="150" swimtime="00:01:48.96" />
                    <SPLIT distance="200" swimtime="00:02:28.21" />
                    <SPLIT distance="250" swimtime="00:03:07.40" />
                    <SPLIT distance="300" swimtime="00:03:46.71" />
                    <SPLIT distance="350" swimtime="00:04:25.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Bessa" birthdate="2003-06-19" gender="M" nation="BRA" license="317841" swrid="5312237" athleteid="2460" externalid="317841">
              <RESULTS>
                <RESULT eventid="1096" points="589" swimtime="00:00:29.75" resultid="2461" heatid="3116" lane="3" entrytime="00:00:29.52" entrycourse="SCM" />
                <RESULT eventid="1320" points="605" reactiontime="+83" swimtime="00:01:05.35" resultid="3300" heatid="3188" lane="4" entrytime="00:01:04.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Antonio Mendes" birthdate="2008-12-04" gender="M" nation="BRA" license="366962" swrid="5196287" athleteid="2513" externalid="366962">
              <RESULTS>
                <RESULT eventid="1096" points="527" swimtime="00:00:30.88" resultid="2514" heatid="3116" lane="2" entrytime="00:00:31.31" entrycourse="SCM" />
                <RESULT eventid="1198" points="320" swimtime="00:20:38.02" resultid="3301" heatid="3150" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:13.58" />
                    <SPLIT distance="150" swimtime="00:01:55.07" />
                    <SPLIT distance="200" swimtime="00:02:36.35" />
                    <SPLIT distance="250" swimtime="00:03:18.57" />
                    <SPLIT distance="300" swimtime="00:03:59.97" />
                    <SPLIT distance="350" swimtime="00:04:41.73" />
                    <SPLIT distance="400" swimtime="00:05:24.21" />
                    <SPLIT distance="450" swimtime="00:06:06.67" />
                    <SPLIT distance="500" swimtime="00:06:48.61" />
                    <SPLIT distance="550" swimtime="00:07:30.24" />
                    <SPLIT distance="600" swimtime="00:08:12.17" />
                    <SPLIT distance="650" swimtime="00:08:54.50" />
                    <SPLIT distance="700" swimtime="00:09:36.79" />
                    <SPLIT distance="750" swimtime="00:10:18.95" />
                    <SPLIT distance="800" swimtime="00:11:01.17" />
                    <SPLIT distance="850" swimtime="00:11:42.82" />
                    <SPLIT distance="900" swimtime="00:12:24.54" />
                    <SPLIT distance="950" swimtime="00:13:06.35" />
                    <SPLIT distance="1000" swimtime="00:13:48.79" />
                    <SPLIT distance="1050" swimtime="00:14:30.87" />
                    <SPLIT distance="1100" swimtime="00:15:12.70" />
                    <SPLIT distance="1150" swimtime="00:15:53.62" />
                    <SPLIT distance="1200" swimtime="00:16:34.66" />
                    <SPLIT distance="1250" swimtime="00:17:15.94" />
                    <SPLIT distance="1300" swimtime="00:17:57.30" />
                    <SPLIT distance="1350" swimtime="00:18:38.97" />
                    <SPLIT distance="1400" swimtime="00:19:20.56" />
                    <SPLIT distance="1450" swimtime="00:20:01.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="545" swimtime="00:01:07.67" resultid="3302" heatid="3188" lane="2" entrytime="00:01:08.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Campelo" birthdate="2011-09-12" gender="M" nation="BRA" license="366963" swrid="5588742" athleteid="2472" externalid="366963">
              <RESULTS>
                <RESULT eventid="1162" points="487" swimtime="00:00:25.61" resultid="2473" heatid="3143" lane="2" entrytime="00:00:25.86" entrycourse="SCM" />
                <RESULT eventid="1140" points="420" reactiontime="+192" swimtime="00:00:29.04" resultid="2474" heatid="3130" lane="2" entrytime="00:00:28.96" entrycourse="SCM" />
                <RESULT eventid="1346" points="474" swimtime="00:00:57.50" resultid="3303" heatid="3203" lane="1" entrytime="00:00:58.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1294" points="394" reactiontime="+77" swimtime="00:00:30.14" resultid="3304" heatid="3178" lane="3" entrytime="00:00:29.89" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolas" lastname="Baldo De França" birthdate="2014-04-21" gender="M" nation="BRA" license="393773" swrid="5507467" athleteid="2649" externalid="393773">
              <RESULTS>
                <RESULT eventid="1151" points="64" swimtime="00:00:50.26" resultid="2650" heatid="3134" lane="2" entrytime="00:00:42.43" entrycourse="SCM" />
                <RESULT eventid="1129" points="76" swimtime="00:00:51.16" resultid="2651" heatid="3127" lane="5" entrytime="00:00:46.86" entrycourse="SCM" />
                <RESULT eventid="1085" points="86" swimtime="00:00:56.43" resultid="2652" heatid="3110" lane="4" entrytime="00:00:56.48" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Yumi Boso" birthdate="2017-11-26" gender="F" nation="BRA" license="421908" athleteid="2778" externalid="421908">
              <RESULTS>
                <RESULT eventid="1276" points="58" swimtime="00:00:30.60" resultid="3305" heatid="3169" lane="5" />
                <RESULT eventid="1228" points="35" swimtime="00:00:34.03" resultid="3306" heatid="3157" lane="4" />
                <RESULT eventid="1302" points="66" swimtime="00:00:32.50" resultid="3307" heatid="3179" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Isabel Henriques" birthdate="2007-09-05" gender="F" nation="BRA" license="414491" swrid="5755356" athleteid="2725" externalid="414491">
              <RESULTS>
                <RESULT eventid="1154" points="206" swimtime="00:00:38.79" resultid="2726" heatid="3137" lane="6" entrytime="00:00:39.65" entrycourse="SCM" />
                <RESULT eventid="1286" points="132" reactiontime="+70" swimtime="00:00:49.58" resultid="3308" heatid="3175" lane="4" entrytime="00:00:48.55" />
                <RESULT eventid="1338" points="174" swimtime="00:01:29.90" resultid="3309" heatid="3196" lane="5" entrytime="00:01:30.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Fernandes Rivadavia" birthdate="2015-11-15" gender="F" nation="BRA" license="393774" swrid="5651342" athleteid="2653" externalid="393774">
              <RESULTS>
                <RESULT eventid="1206" points="217" swimtime="00:01:23.57" resultid="3310" heatid="3152" lane="3" entrytime="00:01:34.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="168" swimtime="00:00:44.13" resultid="3311" heatid="3164" lane="3" entrytime="00:00:51.40" />
                <RESULT eventid="1306" points="167" swimtime="00:00:51.47" resultid="3312" heatid="3182" lane="3" entrytime="00:00:53.96" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio" lastname="Rafael Padial" birthdate="2014-03-07" gender="M" nation="BRA" license="397331" swrid="5641774" athleteid="2665" externalid="397331">
              <RESULTS>
                <RESULT eventid="1151" points="185" swimtime="00:00:35.37" resultid="2666" heatid="3135" lane="5" entrytime="00:00:35.06" entrycourse="SCM" />
                <RESULT eventid="1107" points="144" reactiontime="+80" swimtime="00:00:42.09" resultid="2667" heatid="3120" lane="5" entrytime="00:00:42.10" entrycourse="SCM" />
                <RESULT eventid="1180" points="131" swimtime="00:03:35.76" resultid="3313" heatid="3147" lane="1" entrytime="00:03:26.86" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Munhos Donato" birthdate="2016-07-11" gender="F" nation="BRA" license="421912" athleteid="2794" externalid="421912">
              <RESULTS>
                <RESULT eventid="1254" points="42" swimtime="00:01:09.94" resultid="3314" heatid="3164" lane="2" />
                <RESULT eventid="1280" points="59" reactiontime="+75" swimtime="00:01:04.83" resultid="3315" heatid="3172" lane="6" />
                <RESULT eventid="1332" points="73" swimtime="00:00:54.75" resultid="3316" heatid="3191" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Andrade Silva" birthdate="2016-03-15" gender="M" nation="BRA" license="414852" swrid="5755349" athleteid="2741" externalid="414852">
              <RESULTS>
                <RESULT eventid="1209" points="131" swimtime="00:01:28.16" resultid="3317" heatid="3153" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="106" swimtime="00:01:43.90" resultid="3318" heatid="3160" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1283" points="130" reactiontime="+63" swimtime="00:00:43.55" resultid="3319" heatid="3174" lane="2" entrytime="00:00:49.34" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Beffa Silva" birthdate="2017-02-19" gender="M" nation="BRA" license="421902" athleteid="2754" externalid="421902">
              <RESULTS>
                <RESULT eventid="1230" points="27" swimtime="00:00:32.85" resultid="3320" heatid="3158" lane="5" />
                <RESULT eventid="1304" points="28" swimtime="00:00:37.53" resultid="3321" heatid="3180" lane="4" />
                <RESULT eventid="1330" points="33" swimtime="00:01:02.85" resultid="3322" heatid="3190" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Eduardo Ebiner" birthdate="2013-07-29" gender="M" nation="BRA" license="397371" swrid="5641763" athleteid="2669" externalid="397371">
              <RESULTS>
                <RESULT eventid="1151" status="WDR" swimtime="00:00:00.00" resultid="2670" entrytime="00:00:37.85" entrycourse="SCM" />
                <RESULT eventid="1129" status="WDR" swimtime="00:00:00.00" resultid="2671" entrytime="00:00:43.92" entrycourse="SCM" />
                <RESULT eventid="1085" status="WDR" swimtime="00:00:00.00" resultid="2672" entrytime="00:00:48.17" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Corsine Ferreira" birthdate="2010-03-10" gender="F" nation="BRA" license="353591" swrid="5588608" athleteid="2545" externalid="353591">
              <RESULTS>
                <RESULT eventid="1110" points="330" reactiontime="+63" swimtime="00:01:19.38" resultid="2547" heatid="3122" lane="3" entrytime="00:01:14.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="278" swimtime="00:03:06.64" resultid="3323" heatid="3145" lane="4" entrytime="00:02:51.26" />
                <RESULT eventid="1286" points="309" reactiontime="+68" swimtime="00:00:37.32" resultid="3324" heatid="3176" lane="3" entrytime="00:00:34.06" />
                <RESULT eventid="3234" status="DNS" swimtime="00:00:00.00" resultid="3325" heatid="3754" lane="3" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                    <SPLIT distance="100" swimtime="00:01:22.08" />
                    <SPLIT distance="150" swimtime="00:02:04.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="De Correa" birthdate="2014-12-03" gender="M" nation="BRA" license="403387" swrid="5676286" athleteid="2681" externalid="403387">
              <RESULTS>
                <RESULT eventid="1151" points="168" swimtime="00:00:36.47" resultid="2682" heatid="3134" lane="4" entrytime="00:00:38.51" entrycourse="SCM" />
                <RESULT eventid="1129" points="151" swimtime="00:00:40.79" resultid="2683" heatid="3127" lane="4" entrytime="00:00:42.64" entrycourse="SCM" />
                <RESULT eventid="1107" points="128" swimtime="00:00:43.80" resultid="2684" heatid="3120" lane="6" entrytime="00:00:46.16" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Muniz" birthdate="2012-09-03" gender="M" nation="BRA" license="392106" swrid="5603877" athleteid="2629" externalid="392106">
              <RESULTS>
                <RESULT eventid="1162" points="225" swimtime="00:00:33.14" resultid="2630" heatid="3140" lane="5" entrytime="00:00:34.03" entrycourse="SCM" />
                <RESULT comment="SW 6.4 - Não começou a executar a virada imediatamente após virar para a posição de peito.  (Horário: 9:59), Na volta dos 75m." eventid="1118" reactiontime="+74" status="DSQ" swimtime="00:01:28.86" resultid="2631" heatid="3123" lane="5" entrytime="00:01:45.03" entrycourse="SCM" />
                <RESULT eventid="1346" points="225" swimtime="00:01:13.68" resultid="3326" heatid="3200" lane="1" entrytime="00:01:17.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1294" points="159" reactiontime="+75" swimtime="00:00:40.79" resultid="3327" heatid="3178" lane="6" entrytime="00:00:43.91" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elisa" lastname="Damaziosilva" birthdate="2017-01-26" gender="F" nation="BRA" license="421903" athleteid="2758" externalid="421903">
              <RESULTS>
                <RESULT eventid="1276" points="57" swimtime="00:00:30.68" resultid="3328" heatid="3169" lane="3" />
                <RESULT eventid="1228" points="27" swimtime="00:00:37.12" resultid="3329" heatid="3157" lane="2" />
                <RESULT eventid="1302" points="24" swimtime="00:00:45.24" resultid="3330" heatid="3179" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Rampasi" birthdate="2013-10-16" gender="F" nation="BRA" license="382209" swrid="5603866" athleteid="2609" externalid="382209">
              <RESULTS>
                <RESULT eventid="1060" points="205" swimtime="00:03:06.97" resultid="2610" heatid="3102" lane="1" entrytime="00:03:02.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:02:21.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="206" swimtime="00:00:38.79" resultid="2611" heatid="3132" lane="4" entrytime="00:00:39.77" entrycourse="SCM" />
                <RESULT eventid="1126" points="126" swimtime="00:00:48.59" resultid="2612" heatid="3125" lane="2" entrytime="00:00:48.10" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Amelia Sales" birthdate="2017-07-05" gender="F" nation="BRA" license="421906" athleteid="2770" externalid="421906">
              <RESULTS>
                <RESULT eventid="1276" points="87" swimtime="00:00:26.77" resultid="3331" heatid="3169" lane="1" />
                <RESULT eventid="1228" points="41" swimtime="00:00:32.28" resultid="3332" heatid="3156" lane="4" />
                <RESULT eventid="1328" points="61" swimtime="00:00:58.01" resultid="3333" heatid="3189" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnes" lastname="Sophie Amadei" birthdate="2014-01-10" gender="F" nation="BRA" license="403388" swrid="5676293" athleteid="2685" externalid="403388">
              <RESULTS>
                <RESULT eventid="1060" points="177" swimtime="00:03:16.33" resultid="2686" heatid="3102" lane="6" entrytime="00:03:56.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:02:27.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="190" swimtime="00:00:39.86" resultid="2687" heatid="3132" lane="5" entrytime="00:00:41.94" entrycourse="SCM" />
                <RESULT eventid="1126" points="114" swimtime="00:00:50.15" resultid="2688" heatid="3125" lane="5" entrytime="00:00:51.13" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Campos" birthdate="2013-02-17" gender="M" nation="BRA" license="377262" swrid="5641756" athleteid="2590" externalid="377262">
              <RESULTS>
                <RESULT eventid="1151" points="172" swimtime="00:00:36.19" resultid="2591" heatid="3135" lane="1" entrytime="00:00:35.25" entrycourse="SCM" />
                <RESULT eventid="1107" points="181" reactiontime="+71" swimtime="00:00:39.04" resultid="2592" heatid="3120" lane="3" entrytime="00:00:39.51" entrycourse="SCM" />
                <RESULT eventid="1085" points="140" swimtime="00:00:48.03" resultid="2593" heatid="3111" lane="5" entrytime="00:00:51.31" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietro" lastname="Nabas De Assis" birthdate="2011-07-09" gender="M" nation="BRA" license="366968" swrid="5603878" athleteid="2538" externalid="366968">
              <RESULTS>
                <RESULT eventid="1162" points="313" swimtime="00:00:29.68" resultid="2539" heatid="3141" lane="5" entrytime="00:00:31.03" entrycourse="SCM" />
                <RESULT eventid="1096" points="339" swimtime="00:00:35.77" resultid="2540" heatid="3115" lane="2" entrytime="00:00:34.78" entrycourse="SCM" />
                <RESULT eventid="1346" status="DNS" swimtime="00:00:00.00" resultid="3334" heatid="3199" lane="6" late="yes" />
                <RESULT eventid="1320" status="DNS" swimtime="00:00:00.00" resultid="3335" heatid="3187" lane="3" late="yes" entrytime="00:01:16.01" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tiago" lastname="Ficher Delmont Pais" birthdate="2010-07-15" gender="M" nation="BRA" license="338533" swrid="5588701" athleteid="2468" externalid="338533">
              <RESULTS>
                <RESULT eventid="1180" points="479" swimtime="00:02:20.04" resultid="3336" heatid="3148" lane="3" entrytime="00:02:23.04" />
                <RESULT eventid="1346" points="539" swimtime="00:00:55.09" resultid="3337" heatid="3203" lane="3" entrytime="00:00:55.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" points="429" swimtime="00:05:11.33" resultid="3338" heatid="3155" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                    <SPLIT distance="100" swimtime="00:01:05.44" />
                    <SPLIT distance="150" swimtime="00:01:44.70" />
                    <SPLIT distance="200" swimtime="00:02:24.16" />
                    <SPLIT distance="250" swimtime="00:03:11.59" />
                    <SPLIT distance="300" swimtime="00:04:00.28" />
                    <SPLIT distance="350" swimtime="00:04:36.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniela" lastname="Inoue" birthdate="2008-10-31" gender="F" nation="BRA" license="378348" swrid="5603856" athleteid="2521" externalid="378348">
              <RESULTS>
                <RESULT eventid="1154" points="361" swimtime="00:00:32.19" resultid="2522" heatid="3138" lane="1" entrytime="00:00:31.33" entrycourse="SCM" />
                <RESULT eventid="1110" points="272" reactiontime="+85" swimtime="00:01:24.70" resultid="2523" heatid="3121" lane="3" entrytime="00:01:23.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1338" points="355" swimtime="00:01:10.91" resultid="3339" heatid="3197" lane="3" entrytime="00:01:10.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Bissoli Lucas" birthdate="2017-06-06" gender="M" nation="BRA" license="421907" athleteid="2774" externalid="421907">
              <RESULTS>
                <RESULT eventid="1230" points="17" swimtime="00:00:37.94" resultid="3340" heatid="3158" lane="2" />
                <RESULT eventid="1304" points="31" swimtime="00:00:36.24" resultid="3341" heatid="3180" lane="3" />
                <RESULT eventid="1330" points="18" swimtime="00:01:15.61" resultid="3342" heatid="3190" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduarda" lastname="Pastre" birthdate="2017-09-26" gender="F" nation="BRA" license="421910" athleteid="2786" externalid="421910">
              <RESULTS>
                <RESULT eventid="1276" points="77" swimtime="00:00:27.89" resultid="3343" heatid="3169" lane="6" />
                <RESULT eventid="1228" points="46" swimtime="00:00:31.03" resultid="3344" heatid="3157" lane="1" />
                <RESULT eventid="1328" points="65" swimtime="00:00:56.97" resultid="3345" heatid="3189" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raphael" lastname="Piai Pellegrini" birthdate="2012-03-24" gender="M" nation="BRA" license="377261" swrid="5603894" athleteid="2585" externalid="377261">
              <RESULTS>
                <RESULT eventid="1162" points="358" swimtime="00:00:28.37" resultid="2586" heatid="3142" lane="1" entrytime="00:00:28.98" entrycourse="SCM" />
                <RESULT eventid="1074" points="359" swimtime="00:02:19.69" resultid="2587" heatid="3107" lane="2" entrytime="00:02:24.74" entrycourse="SCM" />
                <RESULT eventid="1346" points="358" swimtime="00:01:03.14" resultid="3346" heatid="3202" lane="6" entrytime="00:01:04.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="242" swimtime="00:01:16.60" resultid="3347" heatid="3168" lane="6" entrytime="00:01:14.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Henrique Goes" birthdate="2008-10-26" gender="M" nation="BRA" license="392105" swrid="5603853" athleteid="2525" externalid="392105">
              <RESULTS>
                <RESULT eventid="1074" points="322" swimtime="00:02:24.91" resultid="2526" heatid="3106" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="100" swimtime="00:01:08.45" />
                    <SPLIT distance="150" swimtime="00:01:46.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="257" swimtime="00:02:52.43" resultid="3348" heatid="3148" lane="1" entrytime="00:02:51.63" />
                <RESULT eventid="1346" points="305" swimtime="00:01:06.56" resultid="3349" heatid="3201" lane="5" entrytime="00:01:07.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="236" swimtime="00:01:17.31" resultid="3350" heatid="3167" lane="3" entrytime="00:01:21.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lara" lastname="Constantino" birthdate="2012-06-02" gender="F" nation="BRA" license="382208" swrid="5420069" athleteid="2604" externalid="382208">
              <RESULTS>
                <RESULT eventid="1154" points="316" swimtime="00:00:33.64" resultid="2605" heatid="3137" lane="3" entrytime="00:00:33.31" entrycourse="SCM" />
                <RESULT eventid="1088" points="318" swimtime="00:00:41.54" resultid="2606" heatid="3112" lane="3" entrytime="00:00:41.26" entrycourse="SCM" />
                <RESULT eventid="1312" points="338" swimtime="00:01:29.44" resultid="3351" heatid="3185" lane="4" entrytime="00:01:31.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1338" points="262" swimtime="00:01:18.52" resultid="3352" heatid="3197" lane="1" entrytime="00:01:17.77" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Catarina" lastname="Wendt Jesus" birthdate="2013-07-09" gender="F" nation="BRA" license="393778" swrid="5641780" athleteid="2661" externalid="393778">
              <RESULTS>
                <RESULT eventid="1060" points="361" swimtime="00:02:34.80" resultid="2662" heatid="3102" lane="3" entrytime="00:02:38.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                    <SPLIT distance="100" swimtime="00:01:16.19" />
                    <SPLIT distance="150" swimtime="00:01:57.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="425" swimtime="00:00:30.48" resultid="2664" heatid="3133" lane="3" entrytime="00:00:31.24" entrycourse="SCM" />
                <RESULT eventid="1170" points="342" swimtime="00:02:54.23" resultid="3353" heatid="3145" lane="5" entrytime="00:02:56.57" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Sunahara Machado" birthdate="2015-03-23" gender="M" nation="BRA" license="421911" athleteid="2790" externalid="421911">
              <RESULTS>
                <RESULT eventid="1283" points="32" swimtime="00:01:09.37" resultid="3354" heatid="3173" lane="2" />
                <RESULT eventid="1309" points="54" swimtime="00:01:05.99" resultid="3355" heatid="3183" lane="3" />
                <RESULT eventid="1335" points="31" swimtime="00:01:03.67" resultid="3356" heatid="3194" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Pedroso Chaim" birthdate="2017-06-14" gender="F" nation="BRA" license="421914" athleteid="2802" externalid="421914">
              <RESULTS>
                <RESULT eventid="1228" points="25" swimtime="00:00:38.11" resultid="3357" heatid="3157" lane="5" />
                <RESULT eventid="1302" points="16" swimtime="00:00:52.28" resultid="3358" heatid="3179" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Marques" birthdate="2015-10-15" gender="F" nation="BRA" license="399738" swrid="5651346" athleteid="2677" externalid="399738">
              <RESULTS>
                <RESULT eventid="1206" points="72" swimtime="00:02:00.69" resultid="3359" heatid="3152" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" points="69" reactiontime="+76" swimtime="00:01:01.40" resultid="3360" heatid="3172" lane="5" entrytime="00:01:08.91" />
                <RESULT eventid="1332" points="70" swimtime="00:00:55.51" resultid="3361" heatid="3193" lane="5" entrytime="00:01:04.05" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Chaim" birthdate="2011-05-29" gender="F" nation="BRA" license="370662" swrid="5409721" athleteid="2553" externalid="370662">
              <RESULTS>
                <RESULT eventid="1154" points="352" swimtime="00:00:32.45" resultid="2554" heatid="3138" lane="6" entrytime="00:00:32.76" entrycourse="SCM" />
                <RESULT eventid="1066" points="342" swimtime="00:02:37.61" resultid="2555" heatid="3105" lane="1" entrytime="00:02:40.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                    <SPLIT distance="100" swimtime="00:01:15.19" />
                    <SPLIT distance="150" swimtime="00:01:56.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="254" reactiontime="+68" swimtime="00:00:39.86" resultid="3362" heatid="3176" lane="5" entrytime="00:00:38.73" />
                <RESULT eventid="1338" points="343" swimtime="00:01:11.72" resultid="3363" heatid="3197" lane="2" entrytime="00:01:12.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Marques Picolo Vinha" birthdate="2010-07-01" gender="M" nation="BRA" license="366990" swrid="5603869" athleteid="2530" externalid="366990">
              <RESULTS>
                <RESULT eventid="1162" points="354" swimtime="00:00:28.48" resultid="2531" heatid="3142" lane="5" entrytime="00:00:28.94" entrycourse="SCM" />
                <RESULT eventid="1346" points="352" swimtime="00:01:03.45" resultid="3364" heatid="3202" lane="5" entrytime="00:01:04.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1246" points="325" swimtime="00:05:08.62" resultid="3365" heatid="3163" lane="2" entrytime="00:05:07.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.06" />
                    <SPLIT distance="100" swimtime="00:01:10.87" />
                    <SPLIT distance="150" swimtime="00:01:50.85" />
                    <SPLIT distance="200" swimtime="00:02:30.65" />
                    <SPLIT distance="250" swimtime="00:03:09.16" />
                    <SPLIT distance="300" swimtime="00:03:49.71" />
                    <SPLIT distance="350" swimtime="00:04:30.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Peroni Passafaro" birthdate="2013-09-17" gender="F" nation="BRA" license="370659" swrid="5603893" athleteid="2567" externalid="370659">
              <RESULTS>
                <RESULT eventid="1126" points="199" swimtime="00:00:41.74" resultid="2569" heatid="3126" lane="2" entrytime="00:00:40.41" entrycourse="SCM" />
                <RESULT eventid="1104" points="259" reactiontime="+72" swimtime="00:00:39.58" resultid="2570" heatid="3117" lane="3" entrytime="00:00:45.15" entrycourse="SCM" />
                <RESULT eventid="1170" points="207" swimtime="00:03:25.79" resultid="3366" heatid="3144" lane="4" entrytime="00:03:30.44" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Batista Sanchez" birthdate="2009-05-22" gender="M" nation="BRA" license="370668" swrid="5255779" athleteid="2481" externalid="370668">
              <RESULTS>
                <RESULT eventid="1096" points="365" swimtime="00:00:34.89" resultid="2482" heatid="3115" lane="3" entrytime="00:00:34.18" entrycourse="SCM" />
                <RESULT eventid="1180" points="360" swimtime="00:02:34.00" resultid="3367" heatid="3148" lane="4" entrytime="00:02:32.12" />
                <RESULT eventid="1320" points="404" swimtime="00:01:14.72" resultid="3368" heatid="3188" lane="5" entrytime="00:01:11.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Allana" lastname="Araujo Oliveira" birthdate="2017-07-25" gender="F" nation="BRA" license="421905" athleteid="2766" externalid="421905">
              <RESULTS>
                <RESULT eventid="1276" points="128" swimtime="00:00:23.54" resultid="3369" heatid="3169" lane="2" />
                <RESULT eventid="1228" points="81" swimtime="00:00:25.80" resultid="3370" heatid="3156" lane="3" />
                <RESULT eventid="1328" points="70" swimtime="00:00:55.40" resultid="3371" heatid="3189" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Dos Reis Monteiro" birthdate="2014-08-05" gender="M" nation="BRA" license="392095" swrid="5697226" athleteid="2617" externalid="392095">
              <RESULTS>
                <RESULT eventid="1151" points="233" swimtime="00:00:32.76" resultid="2618" heatid="3135" lane="3" entrytime="00:00:32.22" entrycourse="SCM" />
                <RESULT eventid="1107" points="169" reactiontime="+82" swimtime="00:00:39.98" resultid="2619" heatid="3120" lane="2" entrytime="00:00:41.41" entrycourse="SCM" />
                <RESULT eventid="1085" points="233" swimtime="00:00:40.52" resultid="2620" heatid="3111" lane="3" entrytime="00:00:40.93" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Otavio Costa" birthdate="2009-01-28" gender="M" nation="BRA" license="370666" swrid="5603881" athleteid="2534" externalid="370666">
              <RESULTS>
                <RESULT eventid="1162" points="294" swimtime="00:00:30.30" resultid="2535" heatid="3141" lane="4" entrytime="00:00:30.80" entrycourse="SCM" />
                <RESULT eventid="1096" points="268" swimtime="00:00:38.66" resultid="2536" heatid="3114" lane="4" entrytime="00:00:39.58" entrycourse="SCM" />
                <RESULT eventid="1246" points="304" swimtime="00:05:15.58" resultid="3372" heatid="3162" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                    <SPLIT distance="100" swimtime="00:01:15.78" />
                    <SPLIT distance="150" swimtime="00:01:56.83" />
                    <SPLIT distance="200" swimtime="00:02:37.14" />
                    <SPLIT distance="250" swimtime="00:03:17.42" />
                    <SPLIT distance="300" swimtime="00:03:58.23" />
                    <SPLIT distance="350" swimtime="00:04:37.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Biason Santana" birthdate="2009-01-21" gender="M" nation="BRA" license="366969" swrid="5317765" athleteid="2517" externalid="366969">
              <RESULTS>
                <RESULT eventid="1140" points="487" swimtime="00:00:27.64" resultid="2518" heatid="3130" lane="4" entrytime="00:00:27.47" entrycourse="SCM" />
                <RESULT eventid="1074" points="407" swimtime="00:02:14.06" resultid="2519" heatid="3106" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.92" />
                    <SPLIT distance="100" swimtime="00:01:04.39" />
                    <SPLIT distance="150" swimtime="00:01:39.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="428" swimtime="00:01:03.36" resultid="3373" heatid="3168" lane="2" entrytime="00:01:02.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Santos Carraro" birthdate="2014-06-04" gender="M" nation="BRA" license="392097" swrid="5603908" athleteid="2621" externalid="392097">
              <RESULTS>
                <RESULT eventid="1151" points="123" swimtime="00:00:40.43" resultid="2622" heatid="3135" lane="6" entrytime="00:00:36.98" entrycourse="SCM" />
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 10:20), Na volta dos 25m." eventid="1129" status="DSQ" swimtime="00:00:43.89" resultid="2623" heatid="3127" lane="2" entrytime="00:00:43.34" entrycourse="SCM" />
                <RESULT eventid="1180" points="114" swimtime="00:03:45.63" resultid="3374" heatid="3146" lane="3" entrytime="00:03:37.77" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aaron" lastname="Michels Dias" birthdate="2017-07-04" gender="M" nation="BRA" license="421909" athleteid="2782" externalid="421909">
              <RESULTS>
                <RESULT eventid="1230" points="45" swimtime="00:00:27.73" resultid="3375" heatid="3158" lane="3" />
                <RESULT eventid="1278" points="61" swimtime="00:00:26.10" resultid="3376" heatid="3170" lane="4" />
                <RESULT eventid="1330" points="48" swimtime="00:00:55.36" resultid="3377" heatid="3190" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juan" lastname="Bernardo Padua" birthdate="2013-07-15" gender="M" nation="BRA" license="392108" swrid="5305422" athleteid="2634" externalid="392108">
              <RESULTS>
                <RESULT eventid="1063" points="207" swimtime="00:02:47.92" resultid="2635" heatid="3103" lane="3" entrytime="00:02:54.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                    <SPLIT distance="100" swimtime="00:01:19.21" />
                    <SPLIT distance="150" swimtime="00:02:06.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1085" points="192" swimtime="00:00:43.24" resultid="2636" heatid="3111" lane="4" entrytime="00:00:43.32" entrycourse="SCM" />
                <RESULT eventid="1180" points="190" swimtime="00:03:10.69" resultid="3378" heatid="3147" lane="2" entrytime="00:03:10.63" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lavinia" lastname="Bossoni" birthdate="2013-11-03" gender="F" nation="BRA" license="377260" swrid="5343093" athleteid="2581" externalid="377260">
              <RESULTS>
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 10:18), Na volta dos 25m." eventid="1126" status="DSQ" swimtime="00:00:48.99" resultid="2582" heatid="3125" lane="3" entrytime="00:00:46.76" entrycourse="SCM" />
                <RESULT eventid="1104" points="203" swimtime="00:00:42.96" resultid="2583" heatid="3118" lane="6" entrytime="00:00:43.53" entrycourse="SCM" />
                <RESULT eventid="1082" points="232" swimtime="00:00:46.16" resultid="2584" heatid="3109" lane="5" entrytime="00:00:50.19" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Quental De Meireles" birthdate="2008-11-20" gender="M" nation="BRA" license="392103" swrid="5603898" athleteid="2543" externalid="392103">
              <RESULTS>
                <RESULT eventid="1268" status="DNS" swimtime="00:00:00.00" resultid="3379" heatid="3168" lane="5" late="yes" entrytime="00:01:07.49" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Pacheco" birthdate="2012-10-03" gender="M" nation="BRA" license="370663" swrid="5603883" athleteid="2571" externalid="370663">
              <RESULTS>
                <RESULT eventid="1162" points="267" swimtime="00:00:31.27" resultid="2572" heatid="3141" lane="6" entrytime="00:00:31.72" entrycourse="SCM" />
                <RESULT eventid="1118" points="209" reactiontime="+64" swimtime="00:01:21.33" resultid="2573" heatid="3123" lane="2" entrytime="00:01:25.93" entrycourse="SCM" />
                <RESULT eventid="1268" points="200" swimtime="00:01:21.70" resultid="3380" heatid="3167" lane="4" entrytime="00:01:23.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 17:46), Na volta dos 25m." eventid="1320" status="DSQ" swimtime="00:01:30.75" resultid="3381" heatid="3186" lane="4" entrytime="00:01:33.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Pastre" birthdate="2014-03-10" gender="F" nation="BRA" license="403760" swrid="5684593" athleteid="2689" externalid="403760">
              <RESULTS>
                <RESULT eventid="1060" points="229" swimtime="00:03:00.20" resultid="2690" heatid="3101" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                    <SPLIT distance="100" swimtime="00:01:26.57" />
                    <SPLIT distance="150" swimtime="00:02:15.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1126" points="187" swimtime="00:00:42.59" resultid="2691" heatid="3126" lane="6" entrytime="00:00:43.88" entrycourse="SCM" />
                <RESULT eventid="1104" points="238" swimtime="00:00:40.72" resultid="2692" heatid="3118" lane="5" entrytime="00:00:40.03" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathan" lastname="Novak Pinho" birthdate="2012-11-14" gender="M" nation="BRA" license="378199" swrid="5603879" athleteid="2599" externalid="378199">
              <RESULTS>
                <RESULT eventid="1118" points="190" reactiontime="+102" swimtime="00:01:24.05" resultid="2600" heatid="3123" lane="4" entrytime="00:01:25.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="232" swimtime="00:02:41.60" resultid="2601" heatid="3106" lane="3" entrytime="00:02:51.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                    <SPLIT distance="100" swimtime="00:01:17.13" />
                    <SPLIT distance="150" swimtime="00:02:00.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1246" points="268" swimtime="00:05:29.01" resultid="3382" heatid="3162" lane="4" entrytime="00:05:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.49" />
                    <SPLIT distance="100" swimtime="00:01:18.47" />
                    <SPLIT distance="150" swimtime="00:02:00.06" />
                    <SPLIT distance="200" swimtime="00:02:42.02" />
                    <SPLIT distance="250" swimtime="00:03:24.68" />
                    <SPLIT distance="300" swimtime="00:04:07.99" />
                    <SPLIT distance="350" swimtime="00:04:48.91" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 6.4 - Não começou a executar a virada imediatamente após virar para a posição de peito.  (Horário: 17:30), Na volta dos 25m." eventid="1294" reactiontime="+101" status="DSQ" swimtime="00:00:37.71" resultid="3383" heatid="3178" lane="5" entrytime="00:00:38.68" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hammon" lastname="Henrique Costa" birthdate="2008-09-19" gender="M" nation="BRA" license="408703" swrid="5726000" athleteid="2720" externalid="408703">
              <RESULTS>
                <RESULT eventid="1162" points="371" swimtime="00:00:28.04" resultid="2721" heatid="3142" lane="3" entrytime="00:00:28.26" entrycourse="SCM" />
                <RESULT eventid="1096" points="356" swimtime="00:00:35.18" resultid="2722" heatid="3115" lane="5" entrytime="00:00:34.79" entrycourse="SCM" />
                <RESULT eventid="1346" points="335" swimtime="00:01:04.50" resultid="3384" heatid="3201" lane="4" entrytime="00:01:04.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="352" swimtime="00:01:18.27" resultid="3385" heatid="3187" lane="2" entrytime="00:01:18.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Cristina Mussolim" birthdate="2015-05-16" gender="F" nation="BRA" license="421913" athleteid="2798" externalid="421913">
              <RESULTS>
                <RESULT eventid="1306" points="75" swimtime="00:01:07.23" resultid="3386" heatid="3181" lane="4" />
                <RESULT eventid="1280" points="63" reactiontime="+101" swimtime="00:01:03.44" resultid="3387" heatid="3171" lane="2" />
                <RESULT eventid="1332" points="93" swimtime="00:00:50.50" resultid="3388" heatid="3192" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Livia" lastname="Rafaela Sita" birthdate="2015-08-10" gender="F" nation="BRA" license="421959" athleteid="2808" externalid="421959">
              <RESULTS>
                <RESULT eventid="1206" points="107" swimtime="00:01:45.71" resultid="3389" heatid="3152" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" points="101" reactiontime="+118" swimtime="00:00:54.05" resultid="3390" heatid="3171" lane="4" />
                <RESULT eventid="1332" points="119" swimtime="00:00:46.61" resultid="3391" heatid="3191" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Izzo Breschiliare" birthdate="2015-09-23" gender="M" nation="BRA" license="407182" swrid="5718669" athleteid="2705" externalid="407182">
              <RESULTS>
                <RESULT eventid="1257" points="50" swimtime="00:00:58.79" resultid="3392" heatid="3165" lane="2" />
                <RESULT eventid="1283" points="59" reactiontime="+76" swimtime="00:00:56.67" resultid="3393" heatid="3173" lane="4" entrytime="00:01:04.74" />
                <RESULT eventid="1335" points="66" swimtime="00:00:49.73" resultid="3394" heatid="3194" lane="4" entrytime="00:01:00.12" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Mochiutti Carneiro" birthdate="2010-04-22" gender="F" nation="BRA" license="370670" swrid="5588817" athleteid="2549" externalid="370670">
              <RESULTS>
                <RESULT eventid="1154" points="389" swimtime="00:00:31.40" resultid="2550" heatid="3138" lane="4" entrytime="00:00:29.36" entrycourse="SCM" />
                <RESULT eventid="1132" points="369" swimtime="00:00:33.98" resultid="2551" heatid="3128" lane="2" entrytime="00:00:31.98" entrycourse="SCM" />
                <RESULT eventid="1066" points="437" swimtime="00:02:25.30" resultid="2552" heatid="3105" lane="4" entrytime="00:02:21.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                    <SPLIT distance="100" swimtime="00:01:09.74" />
                    <SPLIT distance="150" swimtime="00:01:47.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wellington" lastname="De Lima" birthdate="2008-03-01" gender="M" nation="BRA" license="370024" swrid="5470912" athleteid="2477" externalid="370024">
              <RESULTS>
                <RESULT eventid="1162" points="484" swimtime="00:00:25.66" resultid="2478" heatid="3143" lane="5" entrytime="00:00:25.87" entrycourse="SCM" />
                <RESULT eventid="1096" points="441" swimtime="00:00:32.76" resultid="2479" heatid="3116" lane="6" entrytime="00:00:33.99" entrycourse="SCM" />
                <RESULT eventid="1346" points="520" swimtime="00:00:55.75" resultid="3395" heatid="3203" lane="4" entrytime="00:00:56.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Izzo Campos" birthdate="2017-05-29" gender="M" nation="BRA" license="421960" athleteid="2812" externalid="421960">
              <RESULTS>
                <RESULT eventid="1230" points="25" swimtime="00:00:33.33" resultid="3396" heatid="3158" lane="1" />
                <RESULT eventid="1278" points="40" swimtime="00:00:29.99" resultid="3397" heatid="3170" lane="2" />
                <RESULT eventid="1330" points="49" swimtime="00:00:54.74" resultid="3398" heatid="3190" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabrielle" lastname="Borba" birthdate="2014-06-15" gender="F" nation="BRA" license="385705" swrid="5323267" athleteid="2613" externalid="385705">
              <RESULTS>
                <RESULT eventid="1148" points="185" swimtime="00:00:40.19" resultid="2614" heatid="3132" lane="2" entrytime="00:00:41.21" entrycourse="SCM" />
                <RESULT eventid="1126" points="110" swimtime="00:00:50.78" resultid="2615" heatid="3125" lane="4" entrytime="00:00:47.88" entrycourse="SCM" />
                <RESULT eventid="1082" points="170" swimtime="00:00:51.20" resultid="2616" heatid="3109" lane="6" entrytime="00:00:54.15" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Garcia Cavalcante" birthdate="2011-11-21" gender="M" nation="BRA" license="378200" swrid="5603840" athleteid="2489" externalid="378200">
              <RESULTS>
                <RESULT eventid="1096" points="291" swimtime="00:00:37.61" resultid="2490" heatid="3114" lane="3" entrytime="00:00:38.80" entrycourse="SCM" />
                <RESULT comment="SW 6.4 - Não começou a executar a virada imediatamente após virar para a posição de peito.,  Na volta dos 75m (Costas, Medley Individual)." eventid="1180" status="DSQ" swimtime="00:02:50.81" resultid="3399" heatid="3147" lane="3" entrytime="00:03:01.19" />
                <RESULT eventid="1346" points="276" swimtime="00:01:08.86" resultid="3400" heatid="3201" lane="6" entrytime="00:01:09.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="311" swimtime="00:01:21.58" resultid="3401" heatid="3187" lane="1" entrytime="00:01:22.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Guilherme Ortega" birthdate="1999-08-05" gender="M" nation="BRA" license="383118" swrid="5603852" athleteid="2563" externalid="383118">
              <RESULTS>
                <RESULT eventid="1140" points="358" swimtime="00:00:30.61" resultid="2564" heatid="3130" lane="1" entrytime="00:00:30.66" entrycourse="SCM" />
                <RESULT eventid="1180" points="328" swimtime="00:02:38.92" resultid="3402" heatid="3148" lane="2" entrytime="00:02:40.71" />
                <RESULT eventid="1294" points="356" reactiontime="+72" swimtime="00:00:31.19" resultid="3403" heatid="3178" lane="4" entrytime="00:00:30.98" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Passafaro" birthdate="2009-02-01" gender="F" nation="BRA" license="370673" swrid="5603885" athleteid="2504" externalid="370673">
              <RESULTS>
                <RESULT eventid="1154" points="297" swimtime="00:00:34.34" resultid="2505" heatid="3138" lane="5" entrytime="00:00:30.77" entrycourse="SCM" />
                <RESULT eventid="1132" points="336" swimtime="00:00:35.05" resultid="2506" heatid="3128" lane="5" entrytime="00:00:33.10" entrycourse="SCM" />
                <RESULT eventid="1338" points="333" swimtime="00:01:12.45" resultid="3404" heatid="3198" lane="6" entrytime="00:01:09.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Casavechia Carraro" birthdate="2009-07-28" gender="M" nation="BRA" license="368150" swrid="5384752" athleteid="2463" externalid="368150">
              <RESULTS>
                <RESULT eventid="1096" points="415" swimtime="00:00:33.44" resultid="2464" heatid="3116" lane="1" entrytime="00:00:33.54" entrycourse="SCM" />
                <RESULT eventid="1074" points="638" swimtime="00:01:55.38" resultid="2465" heatid="3107" lane="3" entrytime="00:02:00.43" entrycourse="SCM" />
                <RESULT eventid="1246" points="482" swimtime="00:04:30.65" resultid="3405" heatid="3163" lane="3" entrytime="00:04:21.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                    <SPLIT distance="100" swimtime="00:01:02.11" />
                    <SPLIT distance="150" swimtime="00:01:36.12" />
                    <SPLIT distance="200" swimtime="00:02:11.23" />
                    <SPLIT distance="250" swimtime="00:02:46.19" />
                    <SPLIT distance="300" swimtime="00:03:20.64" />
                    <SPLIT distance="350" swimtime="00:03:55.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="504" swimtime="00:01:00.02" resultid="3406" heatid="3168" lane="3" entrytime="00:00:57.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Meneghetti Vidal" birthdate="2015-06-12" gender="M" nation="BRA" license="414851" swrid="5757894" athleteid="2737" externalid="414851">
              <RESULTS>
                <RESULT eventid="1209" points="134" swimtime="00:01:27.60" resultid="3407" heatid="3154" lane="2" entrytime="00:01:35.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="89" swimtime="00:00:48.56" resultid="3408" heatid="3165" lane="4" entrytime="00:00:54.77" />
                <RESULT eventid="1335" points="139" swimtime="00:00:38.86" resultid="3409" heatid="3195" lane="5" entrytime="00:00:42.56" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Otavio Luz" birthdate="2013-07-27" gender="M" nation="BRA" license="392111" swrid="5603882" athleteid="2642" externalid="392111">
              <RESULTS>
                <RESULT eventid="1151" points="227" swimtime="00:00:33.03" resultid="2643" heatid="3135" lane="4" entrytime="00:00:34.34" entrycourse="SCM" />
                <RESULT eventid="1129" points="167" swimtime="00:00:39.49" resultid="2644" heatid="3127" lane="3" entrytime="00:00:38.11" entrycourse="SCM" />
                <RESULT eventid="1107" points="184" reactiontime="+70" swimtime="00:00:38.86" resultid="2645" heatid="3120" lane="4" entrytime="00:00:40.69" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Sanches Ghelere" birthdate="2008-08-06" gender="F" nation="BRA" license="372024" swrid="5603905" athleteid="2508" externalid="372024">
              <RESULTS>
                <RESULT eventid="1154" points="495" swimtime="00:00:28.97" resultid="2509" heatid="3136" lane="2" />
                <RESULT eventid="1132" points="497" swimtime="00:00:30.76" resultid="2510" heatid="3128" lane="4" entrytime="00:00:31.78" entrycourse="SCM" />
                <RESULT eventid="1238" points="477" swimtime="00:04:55.99" resultid="3410" heatid="3161" lane="4" entrytime="00:05:04.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                    <SPLIT distance="100" swimtime="00:01:08.41" />
                    <SPLIT distance="150" swimtime="00:01:45.47" />
                    <SPLIT distance="200" swimtime="00:02:22.61" />
                    <SPLIT distance="250" swimtime="00:02:59.42" />
                    <SPLIT distance="300" swimtime="00:03:35.82" />
                    <SPLIT distance="350" swimtime="00:04:10.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1338" points="515" swimtime="00:01:02.65" resultid="3411" heatid="3198" lane="4" entrytime="00:01:04.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Ghelere" birthdate="2011-04-03" gender="F" nation="BRA" license="368146" swrid="5603843" athleteid="2558" externalid="368146">
              <RESULTS>
                <RESULT eventid="1132" status="SICK" swimtime="00:00:00.00" resultid="2559" entrytime="00:00:36.18" entrycourse="SCM" />
                <RESULT eventid="1110" status="SICK" swimtime="00:00:00.00" resultid="2560" entrytime="00:01:21.65" entrycourse="SCM" />
                <RESULT eventid="1286" status="SICK" swimtime="00:00:00.00" resultid="3412" entrytime="00:00:38.78" />
                <RESULT eventid="1338" status="SICK" swimtime="00:00:00.00" resultid="3413" entrytime="00:01:10.95" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Bassil" birthdate="2015-07-02" gender="M" nation="BRA" license="407178" swrid="5718890" athleteid="2697" externalid="407178">
              <RESULTS>
                <RESULT eventid="1209" points="102" swimtime="00:01:35.93" resultid="3414" heatid="3154" lane="1" entrytime="00:01:47.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1309" points="90" swimtime="00:00:55.50" resultid="3415" heatid="3184" lane="2" entrytime="00:00:56.57" />
                <RESULT eventid="1335" points="103" swimtime="00:00:42.89" resultid="3416" heatid="3195" lane="1" entrytime="00:00:43.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Felipe Sakaguti" birthdate="2007-06-22" gender="M" nation="BRA" license="407187" swrid="5688778" athleteid="2716" externalid="407187">
              <RESULTS>
                <RESULT eventid="1162" points="136" swimtime="00:00:39.16" resultid="2717" heatid="3139" lane="5" entrytime="00:00:42.03" entrycourse="SCM" />
                <RESULT eventid="1346" points="124" swimtime="00:01:29.70" resultid="3417" heatid="3199" lane="4" entrytime="00:01:33.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1294" points="104" reactiontime="+78" swimtime="00:00:46.91" resultid="3418" heatid="3177" lane="4" entrytime="00:00:48.75" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15969" nation="USA" clubid="2821" name="Estados Unidos Da América" shortname="EUA">
          <ATHLETES>
            <ATHLETE firstname="Sophia" lastname="Alanis Whitney" birthdate="2007-07-21" gender="F" nation="USA" license="V397028" swrid="5757088" athleteid="2822" externalid="V397028">
              <RESULTS>
                <RESULT eventid="1154" points="497" swimtime="00:00:28.94" resultid="2823" heatid="3136" lane="4" />
                <RESULT eventid="1132" points="545" swimtime="00:00:29.84" resultid="2824" heatid="3128" lane="3" entrytime="00:00:29.62" entrycourse="SCM" />
                <RESULT eventid="1260" points="556" swimtime="00:01:05.73" resultid="3420" heatid="3166" lane="3" entrytime="00:01:06.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1338" points="501" swimtime="00:01:03.25" resultid="3421" heatid="3198" lane="3" entrytime="00:01:03.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16053" nation="BRA" region="PR" clubid="2827" swrid="93777" name="Fábrica De Nadadores" shortname="Fábrica">
          <ATHLETES>
            <ATHLETE firstname="Eric" lastname="Moreschi" birthdate="2012-08-09" gender="M" nation="BRA" license="385715" swrid="5603876" athleteid="2877" externalid="385715">
              <RESULTS>
                <RESULT eventid="1162" points="245" swimtime="00:00:32.18" resultid="2878" heatid="3140" lane="2" entrytime="00:00:33.29" entrycourse="SCM" />
                <RESULT eventid="1074" points="235" swimtime="00:02:40.92" resultid="2879" heatid="3107" lane="6" entrytime="00:02:48.48" entrycourse="SCM" />
                <RESULT eventid="1246" points="268" swimtime="00:05:29.15" resultid="3422" heatid="3162" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                    <SPLIT distance="100" swimtime="00:01:18.87" />
                    <SPLIT distance="150" swimtime="00:02:00.42" />
                    <SPLIT distance="200" swimtime="00:02:43.44" />
                    <SPLIT distance="250" swimtime="00:03:25.75" />
                    <SPLIT distance="300" swimtime="00:04:07.44" />
                    <SPLIT distance="350" swimtime="00:04:49.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="174" swimtime="00:01:25.53" resultid="3423" heatid="3167" lane="5" entrytime="00:01:31.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marco" lastname="Manzotti Marchi" birthdate="2015-06-26" gender="M" nation="BRA" license="396849" swrid="5641769" athleteid="2936" externalid="396849">
              <RESULTS>
                <RESULT eventid="1209" points="103" swimtime="00:01:35.45" resultid="3424" heatid="3154" lane="5" entrytime="00:01:40.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="101" swimtime="00:00:46.57" resultid="3425" heatid="3165" lane="3" entrytime="00:00:46.68" />
                <RESULT eventid="1335" points="92" swimtime="00:00:44.65" resultid="3426" heatid="3195" lane="6" entrytime="00:00:44.19" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elen" lastname="Torres Gomes" birthdate="2015-10-15" gender="F" nation="BRA" license="396850" swrid="5641777" athleteid="2940" externalid="396850">
              <RESULTS>
                <RESULT eventid="1206" points="122" swimtime="00:01:41.24" resultid="3427" heatid="3152" lane="4" entrytime="00:01:56.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="94" swimtime="00:02:04.07" resultid="3428" heatid="3159" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1306" points="80" swimtime="00:01:05.58" resultid="3429" heatid="3182" lane="4" entrytime="00:01:03.23" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Gevaerd Verssutti Garcia" birthdate="2013-10-15" gender="F" nation="BRA" license="378404" swrid="5588723" athleteid="2915" externalid="378404">
              <RESULTS>
                <RESULT eventid="1060" points="282" swimtime="00:02:48.11" resultid="2916" heatid="3101" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                    <SPLIT distance="100" swimtime="00:01:21.98" />
                    <SPLIT distance="150" swimtime="00:02:06.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1126" points="255" swimtime="00:00:38.40" resultid="2917" heatid="3126" lane="4" entrytime="00:00:38.76" entrycourse="SCM" />
                <RESULT eventid="1104" points="290" swimtime="00:00:38.14" resultid="2918" heatid="3118" lane="2" entrytime="00:00:39.81" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruna" lastname="Scalise Drapzichinski" birthdate="2012-03-07" gender="F" nation="BRA" license="378349" swrid="5603909" athleteid="2843" externalid="378349">
              <RESULTS>
                <RESULT eventid="1154" points="509" swimtime="00:00:28.70" resultid="2845" heatid="3138" lane="2" entrytime="00:00:30.55" entrycourse="SCM" />
                <RESULT eventid="1170" points="378" swimtime="00:02:48.44" resultid="3430" heatid="3145" lane="3" entrytime="00:02:47.79" />
                <RESULT eventid="1312" points="510" swimtime="00:01:18.04" resultid="3431" heatid="3185" lane="3" entrytime="00:01:22.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1338" points="408" swimtime="00:01:07.74" resultid="3432" heatid="3198" lane="1" entrytime="00:01:09.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Braga" birthdate="2010-05-07" gender="M" nation="BRA" license="378345" swrid="5343953" athleteid="2828" externalid="378345">
              <RESULTS>
                <RESULT eventid="1074" points="384" swimtime="00:02:16.63" resultid="2829" heatid="3106" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.44" />
                    <SPLIT distance="100" swimtime="00:01:05.34" />
                    <SPLIT distance="150" swimtime="00:01:41.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="340" swimtime="00:20:12.94" resultid="3433" heatid="3151" lane="2" entrytime="00:21:07.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.64" />
                    <SPLIT distance="100" swimtime="00:01:11.99" />
                    <SPLIT distance="150" swimtime="00:01:50.81" />
                    <SPLIT distance="200" swimtime="00:02:30.83" />
                    <SPLIT distance="250" swimtime="00:03:10.70" />
                    <SPLIT distance="300" swimtime="00:03:51.17" />
                    <SPLIT distance="350" swimtime="00:04:31.72" />
                    <SPLIT distance="400" swimtime="00:05:12.38" />
                    <SPLIT distance="450" swimtime="00:05:52.82" />
                    <SPLIT distance="500" swimtime="00:06:33.36" />
                    <SPLIT distance="550" swimtime="00:07:13.66" />
                    <SPLIT distance="600" swimtime="00:07:54.53" />
                    <SPLIT distance="650" swimtime="00:08:35.27" />
                    <SPLIT distance="700" swimtime="00:09:15.95" />
                    <SPLIT distance="750" swimtime="00:09:56.61" />
                    <SPLIT distance="800" swimtime="00:10:38.11" />
                    <SPLIT distance="850" swimtime="00:11:19.61" />
                    <SPLIT distance="900" swimtime="00:12:00.05" />
                    <SPLIT distance="950" swimtime="00:12:41.41" />
                    <SPLIT distance="1000" swimtime="00:13:22.71" />
                    <SPLIT distance="1050" swimtime="00:14:03.63" />
                    <SPLIT distance="1100" swimtime="00:14:45.36" />
                    <SPLIT distance="1150" swimtime="00:15:26.71" />
                    <SPLIT distance="1200" swimtime="00:16:07.98" />
                    <SPLIT distance="1250" swimtime="00:16:49.28" />
                    <SPLIT distance="1300" swimtime="00:17:31.22" />
                    <SPLIT distance="1350" swimtime="00:18:12.85" />
                    <SPLIT distance="1400" swimtime="00:18:54.13" />
                    <SPLIT distance="1450" swimtime="00:19:34.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" points="370" swimtime="00:05:27.01" resultid="3434" heatid="3155" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                    <SPLIT distance="100" swimtime="00:01:13.04" />
                    <SPLIT distance="150" swimtime="00:01:59.76" />
                    <SPLIT distance="200" swimtime="00:02:46.44" />
                    <SPLIT distance="250" swimtime="00:03:26.74" />
                    <SPLIT distance="300" swimtime="00:04:09.63" />
                    <SPLIT distance="350" swimtime="00:04:49.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="469" reactiontime="+193" swimtime="00:01:11.15" resultid="3435" heatid="3188" lane="1" entrytime="00:01:12.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eloah" lastname="Juvedi Trindade" birthdate="2011-03-05" gender="F" nation="BRA" license="396829" swrid="5641768" athleteid="2931" externalid="396829">
              <RESULTS>
                <RESULT eventid="1154" points="318" reactiontime="+1190" swimtime="00:00:33.56" resultid="2932" heatid="3137" lane="2" entrytime="00:00:33.38" entrycourse="SCM" />
                <RESULT eventid="1190" points="194" swimtime="00:26:08.88" resultid="3436" heatid="3149" lane="2" entrytime="00:24:16.94" />
                <RESULT eventid="1260" points="145" swimtime="00:01:42.79" resultid="3437" heatid="3166" lane="2" entrytime="00:01:46.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="263" swimtime="00:06:00.76" resultid="3438" heatid="3161" lane="6" entrytime="00:06:16.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                    <SPLIT distance="100" swimtime="00:01:25.00" />
                    <SPLIT distance="200" swimtime="00:02:57.96" />
                    <SPLIT distance="250" swimtime="00:03:45.69" />
                    <SPLIT distance="350" swimtime="00:05:18.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theodoro" lastname="Marques Serra" birthdate="2009-11-24" gender="M" nation="BRA" license="370661" swrid="5603870" athleteid="2862" externalid="370661">
              <RESULTS>
                <RESULT eventid="1118" points="387" reactiontime="+66" swimtime="00:01:06.32" resultid="2863" heatid="3124" lane="3" entrytime="00:01:08.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="439" swimtime="00:18:33.88" resultid="3439" heatid="3151" lane="4" entrytime="00:19:42.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                    <SPLIT distance="100" swimtime="00:01:08.33" />
                    <SPLIT distance="150" swimtime="00:01:45.13" />
                    <SPLIT distance="200" swimtime="00:02:22.55" />
                    <SPLIT distance="250" swimtime="00:02:59.75" />
                    <SPLIT distance="300" swimtime="00:03:36.85" />
                    <SPLIT distance="350" swimtime="00:04:13.83" />
                    <SPLIT distance="400" swimtime="00:04:51.31" />
                    <SPLIT distance="450" swimtime="00:05:28.38" />
                    <SPLIT distance="500" swimtime="00:06:05.58" />
                    <SPLIT distance="550" swimtime="00:06:44.11" />
                    <SPLIT distance="600" swimtime="00:07:20.83" />
                    <SPLIT distance="650" swimtime="00:07:57.98" />
                    <SPLIT distance="700" swimtime="00:08:35.79" />
                    <SPLIT distance="750" swimtime="00:09:12.88" />
                    <SPLIT distance="800" swimtime="00:09:51.16" />
                    <SPLIT distance="850" swimtime="00:10:29.40" />
                    <SPLIT distance="900" swimtime="00:11:07.29" />
                    <SPLIT distance="950" swimtime="00:11:44.94" />
                    <SPLIT distance="1000" swimtime="00:12:23.26" />
                    <SPLIT distance="1050" swimtime="00:13:01.17" />
                    <SPLIT distance="1100" swimtime="00:13:38.85" />
                    <SPLIT distance="1150" swimtime="00:14:16.57" />
                    <SPLIT distance="1200" swimtime="00:14:53.84" />
                    <SPLIT distance="1250" swimtime="00:15:31.10" />
                    <SPLIT distance="1300" swimtime="00:16:08.05" />
                    <SPLIT distance="1350" swimtime="00:16:44.98" />
                    <SPLIT distance="1400" swimtime="00:17:22.52" />
                    <SPLIT distance="1450" swimtime="00:17:59.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1346" points="441" swimtime="00:00:58.89" resultid="3440" heatid="3202" lane="4" entrytime="00:01:00.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1246" points="447" swimtime="00:04:37.39" resultid="3441" heatid="3163" lane="4" entrytime="00:04:47.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                    <SPLIT distance="100" swimtime="00:01:04.17" />
                    <SPLIT distance="150" swimtime="00:01:40.05" />
                    <SPLIT distance="200" swimtime="00:02:16.22" />
                    <SPLIT distance="250" swimtime="00:02:52.44" />
                    <SPLIT distance="300" swimtime="00:03:28.06" />
                    <SPLIT distance="350" swimtime="00:04:03.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Dias Hei" birthdate="2016-01-22" gender="F" nation="BRA" license="414653" swrid="5755351" athleteid="2970" externalid="414653">
              <RESULTS>
                <RESULT eventid="1254" points="54" swimtime="00:01:04.12" resultid="3442" heatid="3164" lane="4" />
                <RESULT eventid="1280" points="32" reactiontime="+92" swimtime="00:01:18.97" resultid="3443" heatid="3171" lane="3" />
                <RESULT eventid="1332" points="49" swimtime="00:01:02.43" resultid="3444" heatid="3193" lane="2" entrytime="00:01:03.87" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Berto" birthdate="2008-10-22" gender="M" nation="BRA" license="378342" swrid="5312223" athleteid="2872" externalid="378342">
              <RESULTS>
                <RESULT eventid="1162" points="339" swimtime="00:00:28.91" resultid="2873" heatid="3142" lane="6" entrytime="00:00:30.16" entrycourse="SCM" />
                <RESULT eventid="1096" points="353" swimtime="00:00:35.28" resultid="2874" heatid="3115" lane="1" entrytime="00:00:36.06" entrycourse="SCM" />
                <RESULT eventid="1268" points="225" swimtime="00:01:18.52" resultid="3445" heatid="3167" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="361" swimtime="00:01:17.57" resultid="3446" heatid="3187" lane="5" entrytime="00:01:18.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Laura Oliveira" birthdate="2014-05-19" gender="F" nation="BRA" license="414179" swrid="5336453" athleteid="2969" externalid="414179" />
            <ATHLETE firstname="Sophia" lastname="Schmeiske Ruivo" birthdate="2013-10-21" gender="F" nation="BRA" license="402006" swrid="5661354" athleteid="2944" externalid="402006">
              <RESULTS>
                <RESULT eventid="1148" points="417" swimtime="00:00:30.68" resultid="2946" heatid="3133" lane="4" entrytime="00:00:33.69" entrycourse="SCM" />
                <RESULT eventid="1082" points="369" swimtime="00:00:39.55" resultid="2947" heatid="3109" lane="3" entrytime="00:00:40.68" entrycourse="SCM" />
                <RESULT eventid="1170" points="273" swimtime="00:03:07.71" resultid="3447" heatid="3144" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eloah" lastname="Frasson" birthdate="2012-06-14" gender="F" nation="BRA" license="378338" swrid="5577016" athleteid="2897" externalid="378338">
              <RESULTS>
                <RESULT eventid="1088" points="349" swimtime="00:00:40.29" resultid="2898" heatid="3112" lane="4" entrytime="00:00:42.00" entrycourse="SCM" />
                <RESULT eventid="1190" points="253" swimtime="00:23:54.65" resultid="3448" heatid="3149" lane="1" />
                <RESULT eventid="1312" points="366" reactiontime="+113" swimtime="00:01:27.15" resultid="3449" heatid="3185" lane="2" entrytime="00:01:33.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1338" status="DNS" swimtime="00:00:00.00" resultid="3450" heatid="3196" lane="3" late="yes" entrytime="00:01:18.64" />
                <RESULT eventid="3238" points="300" swimtime="00:03:20.89" resultid="3451" heatid="3532" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.16" />
                    <SPLIT distance="100" swimtime="00:01:36.99" />
                    <SPLIT distance="150" swimtime="00:02:29.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Magalhães Rezende" birthdate="2010-05-29" gender="F" nation="BRA" license="366960" swrid="5588793" athleteid="2867" externalid="366960">
              <RESULTS>
                <RESULT eventid="1066" points="367" swimtime="00:02:34.05" resultid="2868" heatid="3105" lane="5" entrytime="00:02:37.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                    <SPLIT distance="100" swimtime="00:01:12.78" />
                    <SPLIT distance="150" swimtime="00:01:53.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="306" swimtime="00:22:26.65" resultid="3452" heatid="3149" lane="4" entrytime="00:22:31.63" />
                <RESULT eventid="1238" status="DNS" swimtime="00:00:00.00" resultid="3453" heatid="3161" lane="1" late="yes" entrytime="00:05:34.86" />
                <RESULT eventid="1338" status="DNS" swimtime="00:00:00.00" resultid="3454" heatid="3197" lane="4" late="yes" entrytime="00:01:10.40" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Britto" birthdate="2012-10-04" gender="M" nation="BRA" license="378350" swrid="5588566" athleteid="2852" externalid="378350">
              <RESULTS>
                <RESULT eventid="1118" status="DNS" swimtime="00:00:00.00" resultid="2853" heatid="3124" lane="1" entrytime="00:01:15.63" entrycourse="SCM" />
                <RESULT eventid="1074" status="DNS" swimtime="00:00:00.00" resultid="2854" heatid="3107" lane="5" entrytime="00:02:35.57" entrycourse="SCM" />
                <RESULT eventid="1346" status="DNS" swimtime="00:00:00.00" resultid="3455" heatid="3200" lane="4" late="yes" entrytime="00:01:11.31" />
                <RESULT eventid="1220" status="DNS" swimtime="00:00:00.00" resultid="3456" heatid="3155" lane="4" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Dias Rezende" birthdate="2016-03-04" gender="F" nation="BRA" license="406929" swrid="5631410" athleteid="2960" externalid="406929">
              <RESULTS>
                <RESULT eventid="1306" points="46" swimtime="00:01:19.05" resultid="3457" heatid="3181" lane="3" entrytime="00:01:37.96" />
                <RESULT eventid="1332" points="37" swimtime="00:01:08.48" resultid="3458" heatid="3192" lane="4" entrytime="00:01:13.22" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Ognibeni Paupitz" birthdate="2014-08-08" gender="F" nation="BRA" license="406923" swrid="5718889" athleteid="3090" externalid="406923">
              <RESULTS>
                <RESULT eventid="1060" points="121" swimtime="00:03:42.99" resultid="3095" heatid="3101" lane="3" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.51" />
                    <SPLIT distance="100" swimtime="00:01:46.86" />
                    <SPLIT distance="150" swimtime="00:02:47.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1082" points="119" swimtime="00:00:57.63" resultid="3096" heatid="3108" lane="3" late="yes" entrytime="00:00:55.61" entrycourse="SCM" />
                <RESULT eventid="1148" points="129" swimtime="00:00:45.29" resultid="3097" heatid="3132" lane="6" late="yes" entrytime="00:00:43.36" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Voltarelli Souza" birthdate="2014-07-26" gender="M" nation="BRA" license="410202" swrid="5748710" athleteid="2966" externalid="410202">
              <RESULTS>
                <RESULT eventid="1151" status="WDR" swimtime="00:00:00.00" resultid="2967" entrytime="00:00:38.46" entrycourse="SCM" />
                <RESULT eventid="1129" status="WDR" swimtime="00:00:00.00" resultid="2968" entrytime="00:00:44.92" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Miranda Amorim" birthdate="2016-02-06" gender="F" nation="BRA" license="421991" athleteid="2978" externalid="421991">
              <RESULTS>
                <RESULT eventid="1306" points="79" swimtime="00:01:05.90" resultid="3459" heatid="3181" lane="2" />
                <RESULT eventid="1332" points="62" swimtime="00:00:57.91" resultid="3460" heatid="3192" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Rossi" birthdate="2012-05-21" gender="M" nation="BRA" license="378346" swrid="5603901" athleteid="2906" externalid="378346">
              <RESULTS>
                <RESULT eventid="1162" points="270" swimtime="00:00:31.19" resultid="2907" heatid="3141" lane="1" entrytime="00:00:31.54" entrycourse="SCM" />
                <RESULT eventid="1198" points="235" swimtime="00:22:51.61" resultid="3461" heatid="3150" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.94" />
                    <SPLIT distance="100" swimtime="00:01:24.61" />
                    <SPLIT distance="150" swimtime="00:02:10.19" />
                    <SPLIT distance="200" swimtime="00:02:55.17" />
                    <SPLIT distance="250" swimtime="00:03:41.34" />
                    <SPLIT distance="300" swimtime="00:04:27.29" />
                    <SPLIT distance="350" swimtime="00:05:13.27" />
                    <SPLIT distance="400" swimtime="00:06:00.00" />
                    <SPLIT distance="450" swimtime="00:06:46.59" />
                    <SPLIT distance="500" swimtime="00:07:32.33" />
                    <SPLIT distance="550" swimtime="00:08:18.87" />
                    <SPLIT distance="600" swimtime="00:09:05.55" />
                    <SPLIT distance="650" swimtime="00:09:51.82" />
                    <SPLIT distance="700" swimtime="00:10:38.03" />
                    <SPLIT distance="750" swimtime="00:11:24.03" />
                    <SPLIT distance="800" swimtime="00:12:09.54" />
                    <SPLIT distance="850" swimtime="00:12:55.64" />
                    <SPLIT distance="900" swimtime="00:13:40.70" />
                    <SPLIT distance="950" swimtime="00:14:26.47" />
                    <SPLIT distance="1000" swimtime="00:15:12.05" />
                    <SPLIT distance="1050" swimtime="00:15:58.42" />
                    <SPLIT distance="1100" swimtime="00:16:44.41" />
                    <SPLIT distance="1150" swimtime="00:17:30.33" />
                    <SPLIT distance="1200" swimtime="00:18:16.37" />
                    <SPLIT distance="1250" swimtime="00:19:02.44" />
                    <SPLIT distance="1300" swimtime="00:19:49.45" />
                    <SPLIT distance="1350" swimtime="00:20:34.59" />
                    <SPLIT distance="1400" swimtime="00:21:20.83" />
                    <SPLIT distance="1450" swimtime="00:22:06.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1346" status="DNS" swimtime="00:00:00.00" resultid="3462" heatid="3200" lane="3" late="yes" entrytime="00:01:10.38" />
                <RESULT comment="SW 10.2 - Não completou a distância total da prova.  (Horário: 16:35)" eventid="1246" status="DSQ" swimtime="00:00:00.00" resultid="3463" heatid="3162" lane="3" entrytime="00:05:36.77" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Valentina Gonzaga" birthdate="2014-06-28" gender="F" nation="BRA" license="385709" swrid="5603924" athleteid="3089" externalid="385709">
              <RESULTS>
                <RESULT eventid="1082" points="187" swimtime="00:00:49.59" resultid="3098" heatid="3109" lane="1" late="yes" entrytime="00:00:53.76" entrycourse="SCM" />
                <RESULT eventid="1104" points="169" reactiontime="+74" swimtime="00:00:45.63" resultid="3099" heatid="3117" lane="2" late="yes" entrytime="00:00:47.42" entrycourse="SCM" />
                <RESULT eventid="1170" points="162" swimtime="00:03:43.42" resultid="3464" heatid="3144" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Bilemjian Leszczynski" birthdate="2014-02-22" gender="M" nation="BRA" license="406924" swrid="5631285" athleteid="2952" externalid="406924">
              <RESULTS>
                <RESULT eventid="1063" points="126" swimtime="00:03:17.86" resultid="2953" heatid="3103" lane="2" entrytime="00:03:34.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.90" />
                    <SPLIT distance="100" swimtime="00:01:36.99" />
                    <SPLIT distance="150" swimtime="00:02:29.24" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 10:20)" eventid="1129" status="DSQ" swimtime="00:00:55.56" resultid="2954" heatid="3127" lane="6" />
                <RESULT eventid="1085" points="98" swimtime="00:00:54.00" resultid="2955" heatid="3110" lane="2" entrytime="00:00:56.85" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Bagatim" birthdate="2014-05-27" gender="F" nation="BRA" license="378353" swrid="5236649" athleteid="2911" externalid="378353">
              <RESULTS>
                <RESULT eventid="1060" points="260" swimtime="00:02:52.63" resultid="2912" heatid="3101" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.68" />
                    <SPLIT distance="100" swimtime="00:01:21.87" />
                    <SPLIT distance="150" swimtime="00:02:07.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="280" swimtime="00:00:35.03" resultid="2914" heatid="3133" lane="2" entrytime="00:00:34.23" entrycourse="SCM" />
                <RESULT eventid="1170" points="230" swimtime="00:03:18.65" resultid="3465" heatid="3144" lane="3" entrytime="00:03:24.09" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Correa Mendes" birthdate="2015-05-01" gender="M" nation="BRA" license="422089" athleteid="2981" externalid="422089">
              <RESULTS>
                <RESULT eventid="1309" points="84" swimtime="00:00:56.87" resultid="3466" heatid="3183" lane="2" />
                <RESULT eventid="1335" points="71" swimtime="00:00:48.56" resultid="3467" heatid="3194" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="Jacobsen Donati" birthdate="2011-07-14" gender="M" nation="BRA" license="391851" swrid="5615735" athleteid="2882" externalid="391851">
              <RESULTS>
                <RESULT eventid="1118" points="417" reactiontime="+77" swimtime="00:01:04.65" resultid="2883" heatid="3124" lane="4" entrytime="00:01:08.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="303" swimtime="00:21:00.85" resultid="3468" heatid="3150" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:14.51" />
                    <SPLIT distance="150" swimtime="00:01:55.42" />
                    <SPLIT distance="200" swimtime="00:02:36.95" />
                    <SPLIT distance="250" swimtime="00:03:19.19" />
                    <SPLIT distance="300" swimtime="00:04:01.17" />
                    <SPLIT distance="350" swimtime="00:04:43.13" />
                    <SPLIT distance="400" swimtime="00:05:25.42" />
                    <SPLIT distance="450" swimtime="00:06:07.56" />
                    <SPLIT distance="500" swimtime="00:06:50.51" />
                    <SPLIT distance="550" swimtime="00:07:33.21" />
                    <SPLIT distance="600" swimtime="00:08:15.92" />
                    <SPLIT distance="650" swimtime="00:08:59.62" />
                    <SPLIT distance="700" swimtime="00:09:41.86" />
                    <SPLIT distance="750" swimtime="00:10:23.78" />
                    <SPLIT distance="800" swimtime="00:11:06.54" />
                    <SPLIT distance="850" swimtime="00:11:49.07" />
                    <SPLIT distance="900" swimtime="00:12:31.19" />
                    <SPLIT distance="950" swimtime="00:13:14.10" />
                    <SPLIT distance="1000" swimtime="00:13:56.40" />
                    <SPLIT distance="1050" swimtime="00:14:38.67" />
                    <SPLIT distance="1100" swimtime="00:15:21.75" />
                    <SPLIT distance="1150" swimtime="00:16:05.17" />
                    <SPLIT distance="1200" swimtime="00:16:49.36" />
                    <SPLIT distance="1250" swimtime="00:17:31.64" />
                    <SPLIT distance="1300" swimtime="00:18:14.18" />
                    <SPLIT distance="1350" swimtime="00:18:57.54" />
                    <SPLIT distance="1400" swimtime="00:19:40.30" />
                    <SPLIT distance="1450" swimtime="00:20:22.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1346" points="450" swimtime="00:00:58.48" resultid="3469" heatid="3202" lane="2" entrytime="00:01:01.77" />
                <RESULT eventid="1246" points="361" swimtime="00:04:57.95" resultid="3470" heatid="3163" lane="6" entrytime="00:05:34.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                    <SPLIT distance="100" swimtime="00:01:07.80" />
                    <SPLIT distance="150" swimtime="00:01:45.85" />
                    <SPLIT distance="200" swimtime="00:02:24.23" />
                    <SPLIT distance="250" swimtime="00:03:03.68" />
                    <SPLIT distance="300" swimtime="00:03:41.84" />
                    <SPLIT distance="350" swimtime="00:04:21.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andressa" lastname="Zamarian Gouvea" birthdate="2007-09-18" gender="F" nation="BRA" license="318503" swrid="5603929" athleteid="2833" externalid="318503">
              <RESULTS>
                <RESULT eventid="1110" points="347" reactiontime="+70" swimtime="00:01:18.06" resultid="2834" heatid="3122" lane="4" entrytime="00:01:16.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="332" swimtime="00:21:51.01" resultid="3471" heatid="3149" lane="3" entrytime="00:21:13.00" />
                <RESULT eventid="1238" points="420" swimtime="00:05:08.71" resultid="3472" heatid="3161" lane="2" entrytime="00:05:15.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                    <SPLIT distance="100" swimtime="00:01:11.54" />
                    <SPLIT distance="150" swimtime="00:01:50.83" />
                    <SPLIT distance="200" swimtime="00:02:30.34" />
                    <SPLIT distance="250" swimtime="00:03:09.81" />
                    <SPLIT distance="300" swimtime="00:03:49.88" />
                    <SPLIT distance="350" swimtime="00:04:30.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="395" swimtime="00:00:34.41" resultid="3473" heatid="3176" lane="4" entrytime="00:00:34.57" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dante" lastname="Gabriel Rossi" birthdate="2016-01-19" gender="M" nation="BRA" license="406928" swrid="5718627" athleteid="2956" externalid="406928">
              <RESULTS>
                <RESULT eventid="1209" points="70" swimtime="00:01:48.47" resultid="3474" heatid="3153" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1283" points="67" reactiontime="+66" swimtime="00:00:54.19" resultid="3475" heatid="3173" lane="3" entrytime="00:00:55.56" />
                <RESULT eventid="1335" points="82" swimtime="00:00:46.32" resultid="3476" heatid="3194" lane="3" entrytime="00:00:44.61" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Drapzichinski" birthdate="2015-08-21" gender="M" nation="BRA" license="391848" swrid="5603890" athleteid="2927" externalid="391848">
              <RESULTS>
                <RESULT eventid="1209" points="132" swimtime="00:01:27.92" resultid="3477" heatid="3154" lane="4" entrytime="00:01:33.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="131" swimtime="00:01:36.80" resultid="3478" heatid="3160" lane="3" entrytime="00:01:51.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1283" points="120" reactiontime="+87" swimtime="00:00:44.82" resultid="3479" heatid="3174" lane="3" entrytime="00:00:45.94" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kauana" lastname="De Leal" birthdate="2016-02-20" gender="F" nation="BRA" license="417997" athleteid="2974" externalid="417997">
              <RESULTS>
                <RESULT eventid="1232" points="34" swimtime="00:02:53.23" resultid="3480" heatid="3159" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:21.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1306" points="30" swimtime="00:01:30.54" resultid="3481" heatid="3181" lane="1" />
                <RESULT eventid="1332" points="23" swimtime="00:01:19.65" resultid="3482" heatid="3192" lane="3" entrytime="00:01:11.44" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Kenji Yamaguchi" birthdate="2011-08-25" gender="M" nation="BRA" license="385708" swrid="5603862" athleteid="2887" externalid="385708">
              <RESULTS>
                <RESULT eventid="1180" points="313" swimtime="00:02:41.40" resultid="3483" heatid="3148" lane="6" entrytime="00:02:54.66" />
                <RESULT eventid="1198" status="DNS" swimtime="00:00:00.00" resultid="3484" heatid="3151" lane="6" late="yes" entrytime="00:24:55.06" />
                <RESULT eventid="1220" points="300" swimtime="00:05:50.73" resultid="3485" heatid="3155" lane="3" entrytime="00:05:58.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.78" />
                    <SPLIT distance="100" swimtime="00:01:18.03" />
                    <SPLIT distance="150" swimtime="00:02:03.51" />
                    <SPLIT distance="200" swimtime="00:02:49.41" />
                    <SPLIT distance="250" swimtime="00:03:39.35" />
                    <SPLIT distance="300" swimtime="00:04:29.65" />
                    <SPLIT distance="350" swimtime="00:05:11.83" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 10.2 - Não completou a distância total da prova.  (Horário: 16:54)" eventid="1268" status="DSQ" swimtime="00:00:00.00" resultid="3486" heatid="3168" lane="1" entrytime="00:01:12.24" />
                <RESULT eventid="3225" status="DNS" swimtime="00:00:00.00" resultid="3487" heatid="3530" lane="3" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                    <SPLIT distance="100" swimtime="00:01:15.15" />
                    <SPLIT distance="150" swimtime="00:01:57.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Pollettini Canalli" birthdate="2016-08-03" gender="M" nation="BRA" license="422090" athleteid="2984" externalid="422090">
              <RESULTS>
                <RESULT eventid="1209" points="93" swimtime="00:01:38.75" resultid="3488" heatid="3153" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1309" points="69" swimtime="00:01:00.81" resultid="3489" heatid="3183" lane="4" />
                <RESULT eventid="1335" points="87" swimtime="00:00:45.43" resultid="3490" heatid="3194" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Posser" birthdate="2013-02-07" gender="F" nation="BRA" license="378343" swrid="5603896" athleteid="2902" externalid="378343">
              <RESULTS>
                <RESULT eventid="1148" points="231" swimtime="00:00:37.33" resultid="2903" heatid="3133" lane="6" entrytime="00:00:37.17" entrycourse="SCM" />
                <RESULT eventid="1126" points="209" swimtime="00:00:41.08" resultid="2904" heatid="3126" lane="5" entrytime="00:00:41.97" entrycourse="SCM" />
                <RESULT eventid="1104" points="144" reactiontime="+79" swimtime="00:00:48.16" resultid="2905" heatid="3117" lane="5" entrytime="00:00:48.72" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Guinoza" birthdate="2013-01-06" gender="F" nation="BRA" license="392012" swrid="5510698" athleteid="3091" externalid="392012">
              <RESULTS>
                <RESULT eventid="1082" points="233" swimtime="00:00:46.07" resultid="3092" heatid="3109" lane="2" late="yes" entrytime="00:00:48.61" entrycourse="SCM" />
                <RESULT eventid="1126" points="185" swimtime="00:00:42.76" resultid="3093" heatid="3125" lane="1" late="yes" />
                <RESULT eventid="1148" points="253" reactiontime="+1071" swimtime="00:00:36.24" resultid="3094" heatid="3132" lane="3" late="yes" entrytime="00:00:37.98" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Catarina" lastname="Benassi Galvani" birthdate="2015-04-20" gender="F" nation="BRA" license="422153" athleteid="2988" externalid="422153">
              <RESULTS>
                <RESULT eventid="1306" points="67" swimtime="00:01:09.85" resultid="3491" heatid="3181" lane="5" />
                <RESULT eventid="1332" points="97" swimtime="00:00:49.90" resultid="3492" heatid="3191" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Dias Rezende" birthdate="2016-03-04" gender="F" nation="BRA" license="406930" swrid="5685657" athleteid="2963" externalid="406930">
              <RESULTS>
                <RESULT eventid="1306" points="77" swimtime="00:01:06.63" resultid="3493" heatid="3182" lane="1" entrytime="00:01:10.41" />
                <RESULT eventid="1332" points="54" swimtime="00:01:00.32" resultid="3494" heatid="3193" lane="6" entrytime="00:01:10.99" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robsson" lastname="Tows Oliveira" birthdate="2014-03-05" gender="M" nation="BRA" license="392107" swrid="5603922" athleteid="2948" externalid="392107">
              <RESULTS>
                <RESULT eventid="1063" points="159" swimtime="00:03:03.24" resultid="2949" heatid="3103" lane="4" entrytime="00:03:05.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.27" />
                    <SPLIT distance="100" swimtime="00:01:27.20" />
                    <SPLIT distance="150" swimtime="00:02:16.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="183" swimtime="00:00:35.45" resultid="2950" heatid="3134" lane="3" entrytime="00:00:38.03" entrycourse="SCM" />
                <RESULT eventid="1085" points="138" swimtime="00:00:48.23" resultid="2951" heatid="3111" lane="2" entrytime="00:00:48.40" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Tiemi Yamaguchi" birthdate="2013-02-28" gender="F" nation="BRA" license="385707" swrid="5603920" athleteid="2919" externalid="385707">
              <RESULTS>
                <RESULT eventid="1060" points="302" swimtime="00:02:44.40" resultid="2920" heatid="3102" lane="4" entrytime="00:02:49.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.27" />
                    <SPLIT distance="100" swimtime="00:01:19.18" />
                    <SPLIT distance="150" swimtime="00:02:02.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="298" swimtime="00:00:37.77" resultid="2922" heatid="3118" lane="4" entrytime="00:00:38.55" entrycourse="SCM" />
                <RESULT eventid="1170" points="314" swimtime="00:02:59.22" resultid="3495" heatid="3145" lane="1" entrytime="00:02:58.23" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Pazinato" birthdate="2011-01-05" gender="M" nation="BRA" license="368149" swrid="5603889" athleteid="2892" externalid="368149">
              <RESULTS>
                <RESULT eventid="1118" points="288" reactiontime="+75" swimtime="00:01:13.16" resultid="2893" heatid="3124" lane="5" entrytime="00:01:15.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="258" swimtime="00:22:08.64" resultid="3496" heatid="3151" lane="1" entrytime="00:21:52.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                    <SPLIT distance="100" swimtime="00:01:19.31" />
                    <SPLIT distance="150" swimtime="00:02:02.12" />
                    <SPLIT distance="200" swimtime="00:02:44.92" />
                    <SPLIT distance="250" swimtime="00:03:28.72" />
                    <SPLIT distance="300" swimtime="00:04:12.08" />
                    <SPLIT distance="400" swimtime="00:05:39.67" />
                    <SPLIT distance="450" swimtime="00:06:24.11" />
                    <SPLIT distance="500" swimtime="00:07:09.29" />
                    <SPLIT distance="550" swimtime="00:07:54.45" />
                    <SPLIT distance="650" swimtime="00:09:24.59" />
                    <SPLIT distance="700" swimtime="00:10:09.82" />
                    <SPLIT distance="800" swimtime="00:11:41.37" />
                    <SPLIT distance="850" swimtime="00:12:26.76" />
                    <SPLIT distance="900" swimtime="00:13:11.98" />
                    <SPLIT distance="950" swimtime="00:13:57.61" />
                    <SPLIT distance="1000" swimtime="00:14:44.45" />
                    <SPLIT distance="1050" swimtime="00:15:28.56" />
                    <SPLIT distance="1100" swimtime="00:16:15.22" />
                    <SPLIT distance="1450" swimtime="00:21:27.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1346" points="363" swimtime="00:01:02.85" resultid="3497" heatid="3201" lane="3" entrytime="00:01:04.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1246" points="325" swimtime="00:05:08.48" resultid="3498" heatid="3163" lane="1" entrytime="00:05:24.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                    <SPLIT distance="100" swimtime="00:01:11.49" />
                    <SPLIT distance="150" swimtime="00:01:51.06" />
                    <SPLIT distance="200" swimtime="00:02:31.26" />
                    <SPLIT distance="250" swimtime="00:03:11.58" />
                    <SPLIT distance="300" swimtime="00:03:52.82" />
                    <SPLIT distance="350" swimtime="00:04:32.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monique" lastname="Istake" birthdate="2012-04-03" gender="F" nation="BRA" license="372023" swrid="5603857" athleteid="2857" externalid="372023">
              <RESULTS>
                <RESULT eventid="1066" points="364" swimtime="00:02:34.39" resultid="2858" heatid="3104" lane="3" entrytime="00:02:41.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                    <SPLIT distance="100" swimtime="00:01:12.68" />
                    <SPLIT distance="150" swimtime="00:01:55.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="262" swimtime="00:23:38.43" resultid="3499" heatid="3149" lane="5" />
                <RESULT eventid="1260" points="305" swimtime="00:01:20.23" resultid="3500" heatid="3166" lane="4" entrytime="00:01:19.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="367" swimtime="00:01:27.04" resultid="3501" heatid="3185" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Jupi Takaki" birthdate="2013-03-26" gender="F" nation="BRA" license="391845" swrid="5603861" athleteid="2923" externalid="391845">
              <RESULTS>
                <RESULT eventid="1060" points="289" swimtime="00:02:46.74" resultid="2924" heatid="3102" lane="2" entrytime="00:02:49.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                    <SPLIT distance="100" swimtime="00:01:19.72" />
                    <SPLIT distance="150" swimtime="00:02:03.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="289" swimtime="00:00:34.68" resultid="2925" heatid="3133" lane="5" entrytime="00:00:35.74" entrycourse="SCM" />
                <RESULT eventid="1126" points="330" swimtime="00:00:35.27" resultid="2926" heatid="3126" lane="3" entrytime="00:00:36.53" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benicio" lastname="Garcia" birthdate="2011-09-09" gender="M" nation="BRA" license="378347" swrid="5603842" athleteid="2838" externalid="378347">
              <RESULTS>
                <RESULT eventid="1162" points="282" swimtime="00:00:30.72" resultid="2839" heatid="3141" lane="3" entrytime="00:00:30.76" entrycourse="SCM" />
                <RESULT eventid="1198" points="244" swimtime="00:22:33.59" resultid="3502" heatid="3151" lane="5" entrytime="00:21:41.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.77" />
                    <SPLIT distance="100" swimtime="00:01:19.76" />
                    <SPLIT distance="150" swimtime="00:02:02.58" />
                    <SPLIT distance="200" swimtime="00:02:45.97" />
                    <SPLIT distance="250" swimtime="00:03:29.53" />
                    <SPLIT distance="300" swimtime="00:04:12.42" />
                    <SPLIT distance="350" swimtime="00:04:57.18" />
                    <SPLIT distance="400" swimtime="00:05:41.73" />
                    <SPLIT distance="450" swimtime="00:06:27.46" />
                    <SPLIT distance="500" swimtime="00:07:12.48" />
                    <SPLIT distance="550" swimtime="00:07:58.12" />
                    <SPLIT distance="600" swimtime="00:08:44.16" />
                    <SPLIT distance="650" swimtime="00:09:29.39" />
                    <SPLIT distance="700" swimtime="00:10:15.43" />
                    <SPLIT distance="750" swimtime="00:11:02.51" />
                    <SPLIT distance="800" swimtime="00:11:48.29" />
                    <SPLIT distance="850" swimtime="00:12:34.69" />
                    <SPLIT distance="900" swimtime="00:13:21.05" />
                    <SPLIT distance="950" swimtime="00:14:07.96" />
                    <SPLIT distance="1000" swimtime="00:14:54.12" />
                    <SPLIT distance="1050" swimtime="00:15:41.84" />
                    <SPLIT distance="1100" swimtime="00:16:28.83" />
                    <SPLIT distance="1150" swimtime="00:17:17.17" />
                    <SPLIT distance="1200" swimtime="00:18:04.45" />
                    <SPLIT distance="1250" swimtime="00:18:51.60" />
                    <SPLIT distance="1300" swimtime="00:19:38.28" />
                    <SPLIT distance="1350" swimtime="00:20:23.82" />
                    <SPLIT distance="1400" swimtime="00:21:09.04" />
                    <SPLIT distance="1450" swimtime="00:21:52.36" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 16:07), Na volta dos 25m (Borboleta, Medley Individual)." eventid="1220" status="DSQ" swimtime="00:06:28.50" resultid="3503" heatid="3155" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                    <SPLIT distance="100" swimtime="00:01:31.24" />
                    <SPLIT distance="150" swimtime="00:02:19.36" />
                    <SPLIT distance="200" swimtime="00:03:07.56" />
                    <SPLIT distance="250" swimtime="00:04:05.69" />
                    <SPLIT distance="300" swimtime="00:05:03.21" />
                    <SPLIT distance="350" swimtime="00:05:45.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="196" swimtime="00:01:22.17" resultid="3504" heatid="3167" lane="2" entrytime="00:01:28.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabel" lastname="Rezende" birthdate="2013-12-13" gender="F" nation="BRA" license="370657" swrid="5603900" athleteid="2848" externalid="370657">
              <RESULTS>
                <RESULT eventid="1148" points="257" swimtime="00:00:36.03" resultid="2849" heatid="3133" lane="1" entrytime="00:00:36.79" entrycourse="SCM" />
                <RESULT eventid="1126" points="166" reactiontime="+661" swimtime="00:00:44.31" resultid="2850" heatid="3126" lane="1" entrytime="00:00:43.16" entrycourse="SCM" />
                <RESULT eventid="1104" points="229" reactiontime="+72" swimtime="00:00:41.25" resultid="2851" heatid="3117" lane="4" entrytime="00:00:45.88" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15981" nation="BRA" region="PR" clubid="2426" swrid="93783" name="Quinto Nado" shortname="5º Nado">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Fernanda Iossaqui" birthdate="2014-08-01" gender="F" nation="BRA" license="421517" athleteid="2456" externalid="421517">
              <RESULTS>
                <RESULT eventid="1148" points="166" swimtime="00:00:41.65" resultid="2457" heatid="3131" lane="4" />
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 9:23), Na volta dos 25m." eventid="1082" status="DSQ" swimtime="00:00:54.56" resultid="2458" heatid="3108" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benjamin" lastname="Rinaldi Batistao" birthdate="2010-07-13" gender="M" nation="BRA" license="407035" swrid="5737920" athleteid="2451" externalid="407035">
              <RESULTS>
                <RESULT eventid="1162" points="305" swimtime="00:00:29.92" resultid="2452" heatid="3141" lane="2" entrytime="00:00:31.02" entrycourse="SCM" />
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 10:24), Na volta dos 25m." eventid="1140" status="DSQ" swimtime="00:00:33.05" resultid="2453" heatid="3129" lane="3" entrytime="00:00:34.76" entrycourse="SCM" />
                <RESULT eventid="1346" points="316" swimtime="00:01:05.78" resultid="3240" heatid="3201" lane="1" entrytime="00:01:09.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 16:52), Na volta dos 50m." eventid="1268" status="DSQ" swimtime="00:01:22.09" resultid="3241" heatid="3167" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Kikuchi Fujii" birthdate="2007-01-04" gender="M" nation="BRA" license="297805" swrid="5603863" athleteid="2427" externalid="297805">
              <RESULTS>
                <RESULT eventid="1162" points="533" swimtime="00:00:24.86" resultid="2428" heatid="3143" lane="4" entrytime="00:00:25.31" entrycourse="SCM" />
                <RESULT eventid="1096" points="547" swimtime="00:00:30.50" resultid="2429" heatid="3116" lane="4" entrytime="00:00:30.08" entrycourse="SCM" />
                <RESULT eventid="1346" points="536" swimtime="00:00:55.19" resultid="3242" heatid="3203" lane="2" entrytime="00:00:56.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="597" swimtime="00:01:05.64" resultid="3243" heatid="3188" lane="3" entrytime="00:01:03.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco" lastname="Silva Telles" birthdate="2011-07-19" gender="M" nation="BRA" license="377311" swrid="5603911" athleteid="2442" externalid="377311">
              <RESULTS>
                <RESULT eventid="1074" points="295" swimtime="00:02:29.24" resultid="2443" heatid="3106" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                    <SPLIT distance="100" swimtime="00:01:11.53" />
                    <SPLIT distance="150" swimtime="00:01:50.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="257" swimtime="00:02:52.35" resultid="3244" heatid="3147" lane="4" entrytime="00:03:04.06" />
                <RESULT eventid="1246" points="314" swimtime="00:05:12.23" resultid="3245" heatid="3162" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                    <SPLIT distance="100" swimtime="00:01:15.65" />
                    <SPLIT distance="150" swimtime="00:01:56.31" />
                    <SPLIT distance="200" swimtime="00:02:36.72" />
                    <SPLIT distance="250" swimtime="00:03:17.44" />
                    <SPLIT distance="300" swimtime="00:03:57.51" />
                    <SPLIT distance="350" swimtime="00:04:37.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1320" points="281" swimtime="00:01:24.36" resultid="3246" heatid="3186" lane="3" entrytime="00:01:29.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Clara Bobroff" birthdate="2013-02-09" gender="F" nation="BRA" license="391752" swrid="5419807" athleteid="2447" externalid="391752">
              <RESULTS>
                <RESULT eventid="1060" points="276" swimtime="00:02:49.37" resultid="2448" heatid="3102" lane="5" entrytime="00:02:56.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.40" />
                    <SPLIT distance="100" swimtime="00:01:21.96" />
                    <SPLIT distance="150" swimtime="00:02:06.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1082" points="237" swimtime="00:00:45.78" resultid="2450" heatid="3109" lane="4" entrytime="00:00:48.16" entrycourse="SCM" />
                <RESULT eventid="1170" points="211" swimtime="00:03:24.64" resultid="3247" heatid="3144" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Takemura Couto" birthdate="2010-02-08" gender="F" nation="BRA" license="376950" swrid="5603919" athleteid="2437" externalid="376950">
              <RESULTS>
                <RESULT eventid="1154" points="587" swimtime="00:00:27.38" resultid="2438" heatid="3138" lane="3" entrytime="00:00:29.14" entrycourse="SCM" />
                <RESULT eventid="1066" points="560" swimtime="00:02:13.78" resultid="2439" heatid="3105" lane="2" entrytime="00:02:29.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                    <SPLIT distance="100" swimtime="00:01:06.38" />
                    <SPLIT distance="150" swimtime="00:01:40.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="449" reactiontime="+244" swimtime="00:05:02.03" resultid="3248" heatid="3161" lane="5" entrytime="00:05:21.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                    <SPLIT distance="100" swimtime="00:01:10.19" />
                    <SPLIT distance="150" swimtime="00:01:48.13" />
                    <SPLIT distance="200" swimtime="00:02:26.07" />
                    <SPLIT distance="250" swimtime="00:03:05.02" />
                    <SPLIT distance="300" swimtime="00:03:43.33" />
                    <SPLIT distance="350" swimtime="00:04:22.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1338" points="573" swimtime="00:01:00.48" resultid="3249" heatid="3198" lane="2" entrytime="00:01:04.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Poletti Veiga" birthdate="2010-10-01" gender="F" nation="BRA" license="376951" swrid="5603895" athleteid="2432" externalid="376951">
              <RESULTS>
                <RESULT eventid="1110" points="411" reactiontime="+58" swimtime="00:01:13.77" resultid="2433" heatid="3122" lane="2" entrytime="00:01:16.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" points="574" swimtime="00:02:12.66" resultid="2434" heatid="3105" lane="3" entrytime="00:02:18.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.81" />
                    <SPLIT distance="100" swimtime="00:01:06.09" />
                    <SPLIT distance="150" swimtime="00:01:39.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1238" points="533" swimtime="00:04:45.25" resultid="3250" heatid="3161" lane="3" entrytime="00:04:51.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                    <SPLIT distance="100" swimtime="00:01:09.17" />
                    <SPLIT distance="150" swimtime="00:01:45.80" />
                    <SPLIT distance="200" swimtime="00:02:22.83" />
                    <SPLIT distance="250" swimtime="00:02:59.62" />
                    <SPLIT distance="300" swimtime="00:03:35.96" />
                    <SPLIT distance="350" swimtime="00:04:10.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1338" points="490" swimtime="00:01:03.73" resultid="3251" heatid="3198" lane="5" entrytime="00:01:05.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18151" nation="BRA" region="PR" clubid="2816" swrid="95180" name="Clube Uniao Recreativo Palmense" shortname="Clube União">
          <ATHLETES>
            <ATHLETE firstname="Luiza" lastname="Langaro Spaniol" birthdate="2013-06-18" gender="F" nation="BRA" license="406600" swrid="5074027" athleteid="2817" externalid="406600">
              <RESULTS>
                <RESULT eventid="1060" points="411" swimtime="00:02:28.26" resultid="2818" heatid="3101" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                    <SPLIT distance="100" swimtime="00:01:10.70" />
                    <SPLIT distance="150" swimtime="00:01:49.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="363" swimtime="00:00:35.39" resultid="2820" heatid="3118" lane="3" entrytime="00:00:36.64" entrycourse="SCM" />
                <RESULT eventid="1170" points="390" swimtime="00:02:46.72" resultid="3419" heatid="3145" lane="2" entrytime="00:02:55.84" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
