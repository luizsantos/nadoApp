<?xml version="1.0" encoding="UTF-8"?>
<LENEX revisiondate="2024-12-02" created="2025-04-13T16:31:31" version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.81803">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Colombo" name="Troféu Luciano Cabrine (Infantil/Sênior) 2025" course="LCM" deadline="2025-04-05" entrystartdate="2025-03-18" entrytype="INVITATION" hostclub="Santa Mônica Clube de Campo" hostclub.url="https://santamonica.rec.br/" number="39522" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/newInterface/eventos/39522/" startmethod="1" status="OFFICIAL" timing="AUTOMATIC" touchpad="BOTHSIDE" masters="F" withdrawuntil="2025-04-04" state="PR" nation="BRA" hytek.courseorder="L">
      <AGEDATE value="2025-01-01" type="YEAR" />
      <POOL name="Santa Mônica Clube de Campo" lanemax="9" />
      <FACILITY city="Colombo" name="Santa Mônica Clube de Campo" nation="BRA" state="PR" street="Rodovia Régis Bittencourt, KM 6, 5000" street2="Mauá" zip="83413-663" />
      <POINTTABLE pointtableid="3018" name="AQUA Point Scoring" version="2025" />
      <FEES>
        <FEE currency="BRL" type="LATEENTRY.INDIVIDUAL" value="2800" />
        <FEE currency="BRL" type="LATEENTRY.RELAY" value="11200" />
      </FEES>
      <QUALIFY from="2024-03-22" until="2025-03-22" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99252-0598" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99252-0598" street="Avenida do Batel, 1230" street2="Sala 202" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2025-04-11" daytime="08:55" endtime="13:58" number="1" officialmeeting="08:00" status="OFFICIAL" warmupfrom="07:30" warmupuntil="08:30">
          <EVENTS>
            <EVENT eventid="1063" daytime="08:56" gender="F" number="1" order="1" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1064" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8271" />
                    <RANKING order="2" place="2" resultid="8261" />
                    <RANKING order="3" place="3" resultid="8150" />
                    <RANKING order="4" place="4" resultid="8315" />
                    <RANKING order="5" place="5" resultid="9428" />
                    <RANKING order="6" place="6" resultid="8143" />
                    <RANKING order="7" place="7" resultid="9240" />
                    <RANKING order="8" place="8" resultid="8255" />
                    <RANKING order="9" place="9" resultid="7023" />
                    <RANKING order="10" place="10" resultid="8524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8106" />
                    <RANKING order="2" place="2" resultid="8243" />
                    <RANKING order="3" place="3" resultid="8324" />
                    <RANKING order="4" place="4" resultid="8084" />
                    <RANKING order="5" place="5" resultid="6878" />
                    <RANKING order="6" place="6" resultid="9369" />
                    <RANKING order="7" place="7" resultid="7741" />
                    <RANKING order="8" place="8" resultid="7657" />
                    <RANKING order="9" place="9" resultid="6872" />
                    <RANKING order="10" place="10" resultid="8884" />
                    <RANKING order="11" place="11" resultid="7005" />
                    <RANKING order="12" place="12" resultid="9281" />
                    <RANKING order="13" place="-1" resultid="9153" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7594" />
                    <RANKING order="2" place="2" resultid="6565" />
                    <RANKING order="3" place="3" resultid="7987" />
                    <RANKING order="4" place="4" resultid="7098" />
                    <RANKING order="5" place="5" resultid="7219" />
                    <RANKING order="6" place="6" resultid="6994" />
                    <RANKING order="7" place="7" resultid="9307" />
                    <RANKING order="8" place="8" resultid="7768" />
                    <RANKING order="9" place="9" resultid="8979" />
                    <RANKING order="10" place="-1" resultid="9059" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7281" />
                    <RANKING order="2" place="2" resultid="6827" />
                    <RANKING order="3" place="3" resultid="7600" />
                    <RANKING order="4" place="4" resultid="8555" />
                    <RANKING order="5" place="5" resultid="9126" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7921" />
                    <RANKING order="2" place="2" resultid="7398" />
                    <RANKING order="3" place="3" resultid="8965" />
                    <RANKING order="4" place="4" resultid="6959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8679" />
                    <RANKING order="2" place="2" resultid="7333" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10469" daytime="08:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10470" daytime="09:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10471" daytime="09:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10472" daytime="09:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10473" daytime="09:14" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1071" daytime="09:18" gender="M" number="2" order="2" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1072" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8385" />
                    <RANKING order="2" place="2" resultid="7034" />
                    <RANKING order="3" place="3" resultid="7146" />
                    <RANKING order="4" place="4" resultid="8952" />
                    <RANKING order="5" place="5" resultid="8130" />
                    <RANKING order="6" place="6" resultid="8184" />
                    <RANKING order="7" place="7" resultid="8583" />
                    <RANKING order="8" place="8" resultid="8164" />
                    <RANKING order="9" place="9" resultid="8157" />
                    <RANKING order="10" place="10" resultid="8229" />
                    <RANKING order="11" place="11" resultid="7635" />
                    <RANKING order="12" place="12" resultid="8137" />
                    <RANKING order="13" place="13" resultid="7040" />
                    <RANKING order="14" place="14" resultid="9259" />
                    <RANKING order="15" place="15" resultid="7051" />
                    <RANKING order="16" place="-1" resultid="8123" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1073" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7628" />
                    <RANKING order="2" place="2" resultid="8625" />
                    <RANKING order="3" place="3" resultid="8237" />
                    <RANKING order="4" place="4" resultid="9139" />
                    <RANKING order="5" place="5" resultid="7140" />
                    <RANKING order="6" place="6" resultid="8685" />
                    <RANKING order="7" place="7" resultid="8112" />
                    <RANKING order="8" place="8" resultid="7726" />
                    <RANKING order="9" place="9" resultid="8639" />
                    <RANKING order="10" place="10" resultid="8099" />
                    <RANKING order="11" place="11" resultid="8057" />
                    <RANKING order="12" place="12" resultid="9205" />
                    <RANKING order="13" place="13" resultid="9069" />
                    <RANKING order="14" place="-1" resultid="8972" />
                    <RANKING order="15" place="-1" resultid="8711" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1074" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7607" />
                    <RANKING order="2" place="2" resultid="7706" />
                    <RANKING order="3" place="3" resultid="7287" />
                    <RANKING order="4" place="4" resultid="7481" />
                    <RANKING order="5" place="5" resultid="8000" />
                    <RANKING order="6" place="6" resultid="7460" />
                    <RANKING order="7" place="7" resultid="8007" />
                    <RANKING order="8" place="8" resultid="8308" />
                    <RANKING order="9" place="9" resultid="7979" />
                    <RANKING order="10" place="10" resultid="9335" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1075" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7841" />
                    <RANKING order="2" place="2" resultid="7960" />
                    <RANKING order="3" place="3" resultid="7671" />
                    <RANKING order="4" place="4" resultid="8907" />
                    <RANKING order="5" place="5" resultid="8463" />
                    <RANKING order="6" place="6" resultid="7930" />
                    <RANKING order="7" place="-1" resultid="7909" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1076" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7573" />
                    <RANKING order="2" place="2" resultid="7966" />
                    <RANKING order="3" place="-1" resultid="7836" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1077" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7425" />
                    <RANKING order="2" place="2" resultid="8379" />
                    <RANKING order="3" place="3" resultid="8920" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1078" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7419" />
                    <RANKING order="2" place="2" resultid="7561" />
                    <RANKING order="3" place="3" resultid="9593" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10474" daytime="09:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10475" daytime="09:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10476" daytime="09:28" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10477" daytime="09:34" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10478" daytime="09:38" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10479" daytime="09:42" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10480" daytime="09:46" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1079" daytime="09:50" gender="F" number="3" order="3" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1080" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8190" />
                    <RANKING order="2" place="2" resultid="8570" />
                    <RANKING order="3" place="3" resultid="8223" />
                    <RANKING order="4" place="4" resultid="8354" />
                    <RANKING order="5" place="5" resultid="9266" />
                    <RANKING order="6" place="6" resultid="8653" />
                    <RANKING order="7" place="7" resultid="7046" />
                    <RANKING order="8" place="8" resultid="8203" />
                    <RANKING order="9" place="9" resultid="7733" />
                    <RANKING order="10" place="10" resultid="9046" />
                    <RANKING order="11" place="-1" resultid="9211" />
                    <RANKING order="12" place="-1" resultid="6797" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1081" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8064" />
                    <RANKING order="2" place="2" resultid="7691" />
                    <RANKING order="3" place="3" resultid="8070" />
                    <RANKING order="4" place="4" resultid="8331" />
                    <RANKING order="5" place="5" resultid="9132" />
                    <RANKING order="6" place="6" resultid="8078" />
                    <RANKING order="7" place="7" resultid="7761" />
                    <RANKING order="8" place="8" resultid="8513" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7698" />
                    <RANKING order="2" place="2" resultid="7873" />
                    <RANKING order="3" place="3" resultid="8871" />
                    <RANKING order="4" place="4" resultid="9218" />
                    <RANKING order="5" place="5" resultid="8299" />
                    <RANKING order="6" place="6" resultid="9233" />
                    <RANKING order="7" place="7" resultid="8692" />
                    <RANKING order="8" place="8" resultid="6858" />
                    <RANKING order="9" place="9" resultid="8534" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1083" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7935" />
                    <RANKING order="2" place="2" resultid="7879" />
                    <RANKING order="3" place="3" resultid="7310" />
                    <RANKING order="4" place="4" resultid="7822" />
                    <RANKING order="5" place="5" resultid="7940" />
                    <RANKING order="6" place="6" resultid="6837" />
                    <RANKING order="7" place="7" resultid="7446" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1084" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8250" />
                    <RANKING order="2" place="2" resultid="7642" />
                    <RANKING order="3" place="3" resultid="7094" />
                    <RANKING order="4" place="4" resultid="9104" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1085" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8350" />
                    <RANKING order="2" place="2" resultid="7178" />
                    <RANKING order="3" place="3" resultid="9363" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1086" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9531" />
                    <RANKING order="2" place="2" resultid="7580" />
                    <RANKING order="3" place="3" resultid="8878" />
                    <RANKING order="4" place="-1" resultid="8457" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10481" daytime="09:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10482" daytime="09:54" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10483" daytime="10:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10484" daytime="10:04" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10485" daytime="10:08" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10486" daytime="10:12" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1087" daytime="10:18" gender="M" number="4" order="4" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1088" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8285" />
                    <RANKING order="2" place="2" resultid="8177" />
                    <RANKING order="3" place="3" resultid="9191" />
                    <RANKING order="4" place="4" resultid="8210" />
                    <RANKING order="5" place="5" resultid="7754" />
                    <RANKING order="6" place="6" resultid="6931" />
                    <RANKING order="7" place="7" resultid="8170" />
                    <RANKING order="8" place="8" resultid="9329" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1089" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7747" />
                    <RANKING order="2" place="2" resultid="8049" />
                    <RANKING order="3" place="3" resultid="8279" />
                    <RANKING order="4" place="4" resultid="8091" />
                    <RANKING order="5" place="5" resultid="9005" />
                    <RANKING order="6" place="6" resultid="7650" />
                    <RANKING order="7" place="7" resultid="9161" />
                    <RANKING order="8" place="8" resultid="6926" />
                    <RANKING order="9" place="9" resultid="7663" />
                    <RANKING order="10" place="10" resultid="7684" />
                    <RANKING order="11" place="11" resultid="6851" />
                    <RANKING order="12" place="12" resultid="9167" />
                    <RANKING order="13" place="13" resultid="6982" />
                    <RANKING order="14" place="14" resultid="7224" />
                    <RANKING order="15" place="15" resultid="6579" />
                    <RANKING order="16" place="16" resultid="8500" />
                    <RANKING order="17" place="17" resultid="9349" />
                    <RANKING order="18" place="18" resultid="8576" />
                    <RANKING order="19" place="19" resultid="7782" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1090" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8548" />
                    <RANKING order="2" place="2" resultid="9175" />
                    <RANKING order="3" place="3" resultid="8935" />
                    <RANKING order="4" place="4" resultid="9390" />
                    <RANKING order="5" place="5" resultid="7373" />
                    <RANKING order="6" place="6" resultid="7789" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1091" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8913" />
                    <RANKING order="2" place="2" resultid="8394" />
                    <RANKING order="3" place="3" resultid="7299" />
                    <RANKING order="4" place="4" resultid="6914" />
                    <RANKING order="5" place="5" resultid="6976" />
                    <RANKING order="6" place="6" resultid="8475" />
                    <RANKING order="7" place="7" resultid="8782" />
                    <RANKING order="8" place="-1" resultid="7945" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1092" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8267" />
                    <RANKING order="2" place="2" resultid="6946" />
                    <RANKING order="3" place="3" resultid="7678" />
                    <RANKING order="4" place="4" resultid="6920" />
                    <RANKING order="5" place="5" resultid="8959" />
                    <RANKING order="6" place="6" resultid="9053" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1093" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6559" />
                    <RANKING order="2" place="2" resultid="7621" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9512" />
                    <RANKING order="2" place="2" resultid="9564" />
                    <RANKING order="3" place="3" resultid="9599" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10487" daytime="10:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10488" daytime="10:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10489" daytime="10:26" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10490" daytime="10:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10491" daytime="10:34" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10492" daytime="10:38" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1095" daytime="10:42" gender="F" number="5" order="5" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1096" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8590" />
                    <RANKING order="2" place="2" resultid="8569" />
                    <RANKING order="3" place="3" resultid="8736" />
                    <RANKING order="4" place="4" resultid="8652" />
                    <RANKING order="5" place="5" resultid="9427" />
                    <RANKING order="6" place="6" resultid="9239" />
                    <RANKING order="7" place="7" resultid="9045" />
                    <RANKING order="8" place="8" resultid="7157" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1097" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8646" />
                    <RANKING order="2" place="2" resultid="8485" />
                    <RANKING order="3" place="3" resultid="6871" />
                    <RANKING order="4" place="4" resultid="7011" />
                    <RANKING order="5" place="5" resultid="7536" />
                    <RANKING order="6" place="6" resultid="7104" />
                    <RANKING order="7" place="7" resultid="7122" />
                    <RANKING order="8" place="8" resultid="8716" />
                    <RANKING order="9" place="9" resultid="9032" />
                    <RANKING order="10" place="10" resultid="9280" />
                    <RANKING order="11" place="11" resultid="9287" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6572" />
                    <RANKING order="2" place="2" resultid="7195" />
                    <RANKING order="3" place="3" resultid="9181" />
                    <RANKING order="4" place="4" resultid="8985" />
                    <RANKING order="5" place="5" resultid="6999" />
                    <RANKING order="6" place="6" resultid="7872" />
                    <RANKING order="7" place="7" resultid="9299" />
                    <RANKING order="8" place="8" resultid="9586" />
                    <RANKING order="9" place="9" resultid="7593" />
                    <RANKING order="10" place="10" resultid="7923" />
                    <RANKING order="11" place="11" resultid="9232" />
                    <RANKING order="12" place="12" resultid="9306" />
                    <RANKING order="13" place="13" resultid="6866" />
                    <RANKING order="14" place="14" resultid="8978" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1099" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7866" />
                    <RANKING order="2" place="2" resultid="7827" />
                    <RANKING order="3" place="3" resultid="7950" />
                    <RANKING order="4" place="4" resultid="6941" />
                    <RANKING order="5" place="5" resultid="7316" />
                    <RANKING order="6" place="6" resultid="9064" />
                    <RANKING order="7" place="7" resultid="9125" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1100" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7087" />
                    <RANKING order="2" place="2" resultid="7350" />
                    <RANKING order="3" place="3" resultid="8900" />
                    <RANKING order="4" place="4" resultid="9103" />
                    <RANKING order="5" place="5" resultid="7127" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1101" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7177" />
                    <RANKING order="2" place="2" resultid="9083" />
                    <RANKING order="3" place="3" resultid="7565" />
                    <RANKING order="4" place="4" resultid="7332" />
                    <RANKING order="5" place="5" resultid="9362" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7579" />
                    <RANKING order="2" place="2" resultid="9501" />
                    <RANKING order="3" place="3" resultid="9575" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10493" daytime="10:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10494" daytime="10:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10495" daytime="10:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10496" daytime="10:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10497" daytime="10:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10498" daytime="10:52" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1103" daytime="10:54" gender="M" number="6" order="6" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1104" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7028" />
                    <RANKING order="2" place="2" resultid="7322" />
                    <RANKING order="3" place="3" resultid="7017" />
                    <RANKING order="4" place="4" resultid="8216" />
                    <RANKING order="5" place="5" resultid="7356" />
                    <RANKING order="6" place="6" resultid="7171" />
                    <RANKING order="7" place="7" resultid="8618" />
                    <RANKING order="8" place="8" resultid="8659" />
                    <RANKING order="9" place="9" resultid="8742" />
                    <RANKING order="10" place="10" resultid="7501" />
                    <RANKING order="11" place="11" resultid="7251" />
                    <RANKING order="12" place="-1" resultid="7110" />
                    <RANKING order="13" place="-1" resultid="8729" />
                    <RANKING order="14" place="-1" resultid="9225" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1105" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6901" />
                    <RANKING order="2" place="2" resultid="9273" />
                    <RANKING order="3" place="3" resultid="7467" />
                    <RANKING order="4" place="4" resultid="7139" />
                    <RANKING order="5" place="5" resultid="7453" />
                    <RANKING order="6" place="6" resultid="8632" />
                    <RANKING order="7" place="7" resultid="9160" />
                    <RANKING order="8" place="8" resultid="7229" />
                    <RANKING order="9" place="9" resultid="7244" />
                    <RANKING order="10" place="10" resultid="7547" />
                    <RANKING order="11" place="10" resultid="8470" />
                    <RANKING order="12" place="12" resultid="7164" />
                    <RANKING order="13" place="13" resultid="6971" />
                    <RANKING order="14" place="14" resultid="8098" />
                    <RANKING order="15" place="15" resultid="8562" />
                    <RANKING order="16" place="16" resultid="8700" />
                    <RANKING order="17" place="17" resultid="9375" />
                    <RANKING order="18" place="18" resultid="8293" />
                    <RANKING order="19" place="19" resultid="6884" />
                    <RANKING order="20" place="20" resultid="7327" />
                    <RANKING order="21" place="21" resultid="7234" />
                    <RANKING order="22" place="22" resultid="9040" />
                    <RANKING order="23" place="23" resultid="8992" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1106" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9146" />
                    <RANKING order="2" place="2" resultid="8014" />
                    <RANKING order="3" place="3" resultid="8530" />
                    <RANKING order="4" place="4" resultid="9174" />
                    <RANKING order="5" place="5" resultid="9323" />
                    <RANKING order="6" place="6" resultid="9247" />
                    <RANKING order="7" place="7" resultid="7775" />
                    <RANKING order="8" place="8" resultid="9012" />
                    <RANKING order="9" place="9" resultid="7972" />
                    <RANKING order="10" place="10" resultid="8021" />
                    <RANKING order="11" place="11" resultid="9456" />
                    <RANKING order="12" place="12" resultid="9025" />
                    <RANKING order="13" place="13" resultid="9443" />
                    <RANKING order="14" place="14" resultid="7367" />
                    <RANKING order="15" place="15" resultid="9389" />
                    <RANKING order="16" place="-1" resultid="9416" />
                    <RANKING order="17" place="-1" resultid="9422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1107" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6895" />
                    <RANKING order="2" place="2" resultid="8345" />
                    <RANKING order="3" place="3" resultid="7670" />
                    <RANKING order="4" place="4" resultid="8374" />
                    <RANKING order="5" place="5" resultid="6953" />
                    <RANKING order="6" place="6" resultid="8772" />
                    <RANKING order="7" place="7" resultid="8605" />
                    <RANKING order="8" place="8" resultid="9292" />
                    <RANKING order="9" place="9" resultid="7304" />
                    <RANKING order="10" place="10" resultid="7955" />
                    <RANKING order="11" place="11" resultid="9449" />
                    <RANKING order="12" place="-1" resultid="7847" />
                    <RANKING order="13" place="-1" resultid="8491" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1108" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7572" />
                    <RANKING order="2" place="2" resultid="9397" />
                    <RANKING order="3" place="3" resultid="9110" />
                    <RANKING order="4" place="4" resultid="9090" />
                    <RANKING order="5" place="5" resultid="7411" />
                    <RANKING order="6" place="6" resultid="6907" />
                    <RANKING order="7" place="7" resultid="6988" />
                    <RANKING order="8" place="8" resultid="7344" />
                    <RANKING order="9" place="9" resultid="7384" />
                    <RANKING order="10" place="10" resultid="9052" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1109" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6558" />
                    <RANKING order="2" place="2" resultid="8891" />
                    <RANKING order="3" place="3" resultid="6935" />
                    <RANKING order="4" place="4" resultid="8672" />
                    <RANKING order="5" place="5" resultid="7530" />
                    <RANKING order="6" place="6" resultid="9314" />
                    <RANKING order="7" place="7" resultid="8941" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1110" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7200" />
                    <RANKING order="2" place="2" resultid="7418" />
                    <RANKING order="3" place="3" resultid="7205" />
                    <RANKING order="4" place="4" resultid="9519" />
                    <RANKING order="5" place="5" resultid="9544" />
                    <RANKING order="6" place="6" resultid="9550" />
                    <RANKING order="7" place="7" resultid="9598" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10499" daytime="10:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10500" daytime="10:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10501" daytime="10:58" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10502" daytime="11:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10503" daytime="11:02" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10504" daytime="11:04" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10505" daytime="11:04" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10506" daytime="11:06" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10507" daytime="11:08" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10508" daytime="11:10" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1111" daytime="11:22" gender="X" number="7" order="8" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1112" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8433" />
                    <RANKING order="2" place="2" resultid="8452" />
                    <RANKING order="3" place="3" resultid="8755" />
                    <RANKING order="4" place="4" resultid="7077" />
                    <RANKING order="5" place="5" resultid="9484" />
                    <RANKING order="6" place="6" resultid="9493" />
                    <RANKING order="7" place="7" resultid="8759" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10509" daytime="11:22" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1113" daytime="11:28" gender="X" number="8" order="9" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1114" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8432" />
                    <RANKING order="2" place="2" resultid="7816" />
                    <RANKING order="3" place="3" resultid="8451" />
                    <RANKING order="4" place="4" resultid="9483" />
                    <RANKING order="5" place="5" resultid="8754" />
                    <RANKING order="6" place="6" resultid="7800" />
                    <RANKING order="7" place="7" resultid="7076" />
                    <RANKING order="8" place="8" resultid="6891" />
                    <RANKING order="9" place="-1" resultid="9492" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10510" daytime="11:28" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1115" daytime="11:36" gender="F" number="9" order="10" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1116" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8197" />
                    <RANKING order="2" place="2" resultid="8222" />
                    <RANKING order="3" place="3" resultid="9018" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1117" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8077" />
                    <RANKING order="2" place="2" resultid="8063" />
                    <RANKING order="3" place="3" resultid="8105" />
                    <RANKING order="4" place="4" resultid="7656" />
                    <RANKING order="5" place="5" resultid="7740" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1118" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8927" />
                    <RANKING order="2" place="2" resultid="7494" />
                    <RANKING order="3" place="3" resultid="7986" />
                    <RANKING order="4" place="4" resultid="8611" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1119" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7860" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1120" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8400" />
                    <RANKING order="2" place="2" resultid="8964" />
                    <RANKING order="3" place="3" resultid="8899" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1121" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8678" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1122" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8322" />
                    <RANKING order="2" place="2" resultid="8361" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10511" daytime="11:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10512" daytime="11:58" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1123" daytime="12:20" gender="M" number="10" order="11" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1124" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8163" />
                    <RANKING order="2" place="2" resultid="7719" />
                    <RANKING order="3" place="3" resultid="8183" />
                    <RANKING order="4" place="4" resultid="8136" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1125" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8236" />
                    <RANKING order="2" place="2" resultid="7649" />
                    <RANKING order="3" place="3" resultid="8035" />
                    <RANKING order="4" place="4" resultid="8971" />
                    <RANKING order="5" place="5" resultid="9198" />
                    <RANKING order="6" place="6" resultid="8056" />
                    <RANKING order="7" place="7" resultid="9004" />
                    <RANKING order="8" place="8" resultid="8278" />
                    <RANKING order="9" place="9" resultid="8367" />
                    <RANKING order="10" place="10" resultid="9039" />
                    <RANKING order="11" place="-1" resultid="8042" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7902" />
                    <RANKING order="2" place="2" resultid="8028" />
                    <RANKING order="3" place="3" resultid="7705" />
                    <RANKING order="4" place="4" resultid="8934" />
                    <RANKING order="5" place="5" resultid="9246" />
                    <RANKING order="6" place="6" resultid="8946" />
                    <RANKING order="7" place="7" resultid="7614" />
                    <RANKING order="8" place="8" resultid="9011" />
                    <RANKING order="9" place="-1" resultid="7914" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1127" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8906" />
                    <RANKING order="2" place="2" resultid="7885" />
                    <RANKING order="3" place="3" resultid="7586" />
                    <RANKING order="4" place="4" resultid="8604" />
                    <RANKING order="5" place="5" resultid="6842" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8119" />
                    <RANKING order="2" place="2" resultid="7432" />
                    <RANKING order="3" place="3" resultid="7712" />
                    <RANKING order="4" place="4" resultid="7677" />
                    <RANKING order="5" place="5" resultid="9396" />
                    <RANKING order="6" place="6" resultid="8509" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1129" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7893" />
                    <RANKING order="2" place="2" resultid="9313" />
                    <RANKING order="3" place="3" resultid="7439" />
                    <RANKING order="4" place="4" resultid="8671" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1130" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7560" />
                    <RANKING order="2" place="2" resultid="9382" />
                    <RANKING order="3" place="3" resultid="9563" />
                    <RANKING order="4" place="4" resultid="9556" />
                    <RANKING order="5" place="5" resultid="9592" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10513" daytime="12:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10514" daytime="12:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10515" daytime="12:42" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10516" daytime="12:54" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10517" daytime="13:06" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2025-04-11" daytime="16:25" endtime="20:22" number="2" officialmeeting="15:00" status="OFFICIAL" warmupfrom="14:30" warmupuntil="15:30">
          <EVENTS>
            <EVENT eventid="1131" daytime="16:26" gender="F" number="11" order="1" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1132" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8224" />
                    <RANKING order="2" place="2" resultid="8198" />
                    <RANKING order="3" place="3" resultid="8205" />
                    <RANKING order="4" place="4" resultid="7735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1133" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8065" />
                    <RANKING order="2" place="2" resultid="7693" />
                    <RANKING order="3" place="3" resultid="7763" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1134" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7699" />
                    <RANKING order="2" place="2" resultid="8873" />
                    <RANKING order="3" place="3" resultid="8928" />
                    <RANKING order="4" place="4" resultid="7769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1135" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7601" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1136" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7399" />
                    <RANKING order="2" place="2" resultid="8902" />
                    <RANKING order="3" place="-1" resultid="7644" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1137" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8680" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1138" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10518" daytime="16:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10519" daytime="16:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10520" daytime="16:40" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1139" daytime="16:48" gender="M" number="12" order="2" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1140" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7035" />
                    <RANKING order="2" place="2" resultid="7637" />
                    <RANKING order="3" place="3" resultid="8584" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1141" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7651" />
                    <RANKING order="2" place="2" resultid="8113" />
                    <RANKING order="3" place="3" resultid="7728" />
                    <RANKING order="4" place="4" resultid="7665" />
                    <RANKING order="5" place="5" resultid="7749" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1142" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7609" />
                    <RANKING order="2" place="2" resultid="8008" />
                    <RANKING order="3" place="3" resultid="7289" />
                    <RANKING order="4" place="4" resultid="7707" />
                    <RANKING order="5" place="5" resultid="7777" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1143" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8908" />
                    <RANKING order="2" place="2" resultid="7673" />
                    <RANKING order="3" place="3" resultid="7588" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1144" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7574" />
                    <RANKING order="2" place="2" resultid="7433" />
                    <RANKING order="3" place="3" resultid="7679" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1145" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7427" />
                    <RANKING order="2" place="-1" resultid="7623" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1146" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9557" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10521" daytime="16:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10522" daytime="16:54" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10523" daytime="17:02" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1147" daytime="17:08" gender="F" number="13" order="3" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1148" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8151" />
                    <RANKING order="2" place="2" resultid="8144" />
                    <RANKING order="3" place="3" resultid="8262" />
                    <RANKING order="4" place="4" resultid="8355" />
                    <RANKING order="5" place="5" resultid="9241" />
                    <RANKING order="6" place="6" resultid="8572" />
                    <RANKING order="7" place="7" resultid="8204" />
                    <RANKING order="8" place="8" resultid="8737" />
                    <RANKING order="9" place="9" resultid="8316" />
                    <RANKING order="10" place="10" resultid="9429" />
                    <RANKING order="11" place="11" resultid="7133" />
                    <RANKING order="12" place="12" resultid="8256" />
                    <RANKING order="13" place="13" resultid="9604" />
                    <RANKING order="14" place="14" resultid="7024" />
                    <RANKING order="15" place="15" resultid="8191" />
                    <RANKING order="16" place="16" resultid="9047" />
                    <RANKING order="17" place="17" resultid="9019" />
                    <RANKING order="18" place="18" resultid="8789" />
                    <RANKING order="19" place="19" resultid="9213" />
                    <RANKING order="20" place="20" resultid="7159" />
                    <RANKING order="21" place="21" resultid="7362" />
                    <RANKING order="22" place="22" resultid="8525" />
                    <RANKING order="23" place="23" resultid="8666" />
                    <RANKING order="24" place="24" resultid="9411" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1149" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6879" />
                    <RANKING order="2" place="2" resultid="8107" />
                    <RANKING order="3" place="3" resultid="8648" />
                    <RANKING order="4" place="4" resultid="8079" />
                    <RANKING order="5" place="5" resultid="8085" />
                    <RANKING order="6" place="6" resultid="7742" />
                    <RANKING order="7" place="7" resultid="8486" />
                    <RANKING order="8" place="8" resultid="8244" />
                    <RANKING order="9" place="9" resultid="8598" />
                    <RANKING order="10" place="10" resultid="8325" />
                    <RANKING order="11" place="11" resultid="9370" />
                    <RANKING order="12" place="12" resultid="7658" />
                    <RANKING order="13" place="13" resultid="8333" />
                    <RANKING order="14" place="14" resultid="6873" />
                    <RANKING order="15" place="15" resultid="7006" />
                    <RANKING order="16" place="16" resultid="9134" />
                    <RANKING order="17" place="17" resultid="8072" />
                    <RANKING order="18" place="18" resultid="7012" />
                    <RANKING order="19" place="19" resultid="7489" />
                    <RANKING order="20" place="20" resultid="8885" />
                    <RANKING order="21" place="21" resultid="9282" />
                    <RANKING order="22" place="22" resultid="7124" />
                    <RANKING order="23" place="23" resultid="8718" />
                    <RANKING order="24" place="24" resultid="9404" />
                    <RANKING order="25" place="25" resultid="8403" />
                    <RANKING order="26" place="26" resultid="6587" />
                    <RANKING order="27" place="27" resultid="9033" />
                    <RANKING order="28" place="28" resultid="9288" />
                    <RANKING order="29" place="29" resultid="9357" />
                    <RANKING order="30" place="-1" resultid="9154" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6573" />
                    <RANKING order="2" place="2" resultid="6566" />
                    <RANKING order="3" place="3" resultid="7925" />
                    <RANKING order="4" place="4" resultid="7874" />
                    <RANKING order="5" place="5" resultid="7000" />
                    <RANKING order="6" place="6" resultid="7988" />
                    <RANKING order="7" place="7" resultid="9183" />
                    <RANKING order="8" place="8" resultid="9300" />
                    <RANKING order="9" place="9" resultid="7099" />
                    <RANKING order="10" place="10" resultid="7993" />
                    <RANKING order="11" place="11" resultid="7554" />
                    <RANKING order="12" place="12" resultid="9587" />
                    <RANKING order="13" place="13" resultid="8612" />
                    <RANKING order="14" place="14" resultid="7081" />
                    <RANKING order="15" place="15" resultid="8694" />
                    <RANKING order="16" place="16" resultid="7595" />
                    <RANKING order="17" place="17" resultid="9308" />
                    <RANKING order="18" place="18" resultid="7495" />
                    <RANKING order="19" place="19" resultid="6862" />
                    <RANKING order="20" place="20" resultid="6860" />
                    <RANKING order="21" place="21" resultid="6867" />
                    <RANKING order="22" place="22" resultid="9060" />
                    <RANKING order="23" place="23" resultid="8799" />
                    <RANKING order="24" place="24" resultid="8301" />
                    <RANKING order="25" place="25" resultid="7152" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1151" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7828" />
                    <RANKING order="2" place="2" resultid="7861" />
                    <RANKING order="3" place="3" resultid="6828" />
                    <RANKING order="4" place="4" resultid="7951" />
                    <RANKING order="5" place="5" resultid="7282" />
                    <RANKING order="6" place="6" resultid="7318" />
                    <RANKING order="7" place="7" resultid="7215" />
                    <RANKING order="8" place="8" resultid="7524" />
                    <RANKING order="9" place="9" resultid="7448" />
                    <RANKING order="10" place="10" resultid="9127" />
                    <RANKING order="11" place="11" resultid="6942" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1152" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7088" />
                    <RANKING order="2" place="2" resultid="8998" />
                    <RANKING order="3" place="3" resultid="7351" />
                    <RANKING order="4" place="4" resultid="7210" />
                    <RANKING order="5" place="5" resultid="9106" />
                    <RANKING order="6" place="6" resultid="6960" />
                    <RANKING order="7" place="7" resultid="7128" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1153" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9084" />
                    <RANKING order="2" place="2" resultid="7334" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1154" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9526" />
                    <RANKING order="2" place="2" resultid="9576" />
                    <RANKING order="3" place="3" resultid="9503" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10524" daytime="17:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10525" daytime="17:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10526" daytime="17:14" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10527" daytime="17:16" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10528" daytime="17:18" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10529" daytime="17:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10530" daytime="17:22" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10531" daytime="17:24" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10532" daytime="17:26" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10533" daytime="17:28" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="10534" daytime="17:30" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1155" daytime="17:34" gender="M" number="14" order="4" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1156" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7509" />
                    <RANKING order="2" place="2" resultid="8386" />
                    <RANKING order="3" place="3" resultid="7029" />
                    <RANKING order="4" place="4" resultid="8165" />
                    <RANKING order="5" place="5" resultid="7147" />
                    <RANKING order="6" place="6" resultid="8178" />
                    <RANKING order="7" place="7" resultid="8131" />
                    <RANKING order="8" place="7" resultid="8286" />
                    <RANKING order="9" place="9" resultid="7357" />
                    <RANKING order="10" place="10" resultid="9193" />
                    <RANKING order="11" place="11" resultid="8211" />
                    <RANKING order="12" place="12" resultid="9342" />
                    <RANKING order="13" place="13" resultid="7323" />
                    <RANKING order="14" place="14" resultid="8185" />
                    <RANKING order="15" place="15" resultid="8158" />
                    <RANKING order="16" place="16" resultid="8953" />
                    <RANKING order="17" place="17" resultid="7111" />
                    <RANKING order="18" place="18" resultid="7019" />
                    <RANKING order="19" place="19" resultid="7172" />
                    <RANKING order="20" place="20" resultid="8661" />
                    <RANKING order="21" place="21" resultid="7041" />
                    <RANKING order="22" place="22" resultid="8724" />
                    <RANKING order="23" place="23" resultid="7052" />
                    <RANKING order="24" place="24" resultid="8743" />
                    <RANKING order="25" place="25" resultid="8231" />
                    <RANKING order="26" place="26" resultid="8481" />
                    <RANKING order="27" place="27" resultid="7253" />
                    <RANKING order="28" place="28" resultid="7636" />
                    <RANKING order="29" place="29" resultid="9260" />
                    <RANKING order="30" place="30" resultid="7380" />
                    <RANKING order="31" place="31" resultid="7117" />
                    <RANKING order="32" place="32" resultid="7503" />
                    <RANKING order="33" place="33" resultid="8171" />
                    <RANKING order="34" place="34" resultid="9253" />
                    <RANKING order="35" place="35" resultid="9331" />
                    <RANKING order="36" place="36" resultid="9435" />
                    <RANKING order="37" place="37" resultid="8762" />
                    <RANKING order="38" place="38" resultid="8814" />
                    <RANKING order="39" place="39" resultid="8819" />
                    <RANKING order="40" place="-1" resultid="8730" />
                    <RANKING order="41" place="-1" resultid="9226" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1157" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8238" />
                    <RANKING order="2" place="2" resultid="6902" />
                    <RANKING order="3" place="3" resultid="8050" />
                    <RANKING order="4" place="4" resultid="8093" />
                    <RANKING order="5" place="5" resultid="7141" />
                    <RANKING order="6" place="6" resultid="8036" />
                    <RANKING order="7" place="7" resultid="7455" />
                    <RANKING order="8" place="8" resultid="9169" />
                    <RANKING order="9" place="9" resultid="9206" />
                    <RANKING order="10" place="10" resultid="7542" />
                    <RANKING order="11" place="11" resultid="8640" />
                    <RANKING order="12" place="12" resultid="7727" />
                    <RANKING order="13" place="13" resultid="6853" />
                    <RANKING order="14" place="14" resultid="7230" />
                    <RANKING order="15" place="15" resultid="8368" />
                    <RANKING order="16" place="16" resultid="8471" />
                    <RANKING order="17" place="17" resultid="7748" />
                    <RANKING order="18" place="18" resultid="8712" />
                    <RANKING order="19" place="19" resultid="8973" />
                    <RANKING order="20" place="20" resultid="7062" />
                    <RANKING order="21" place="21" resultid="8295" />
                    <RANKING order="22" place="22" resultid="7548" />
                    <RANKING order="23" place="23" resultid="7328" />
                    <RANKING order="24" place="23" resultid="8100" />
                    <RANKING order="25" place="25" resultid="6581" />
                    <RANKING order="26" place="26" resultid="8058" />
                    <RANKING order="27" place="27" resultid="7239" />
                    <RANKING order="28" place="28" resultid="7246" />
                    <RANKING order="29" place="29" resultid="6972" />
                    <RANKING order="30" place="30" resultid="7166" />
                    <RANKING order="31" place="31" resultid="9041" />
                    <RANKING order="32" place="32" resultid="6886" />
                    <RANKING order="33" place="33" resultid="7475" />
                    <RANKING order="34" place="34" resultid="7784" />
                    <RANKING order="35" place="35" resultid="9377" />
                    <RANKING order="36" place="36" resultid="7235" />
                    <RANKING order="37" place="37" resultid="9351" />
                    <RANKING order="38" place="38" resultid="8578" />
                    <RANKING order="39" place="39" resultid="9071" />
                    <RANKING order="40" place="40" resultid="8809" />
                    <RANKING order="41" place="41" resultid="8707" />
                    <RANKING order="42" place="42" resultid="8768" />
                    <RANKING order="43" place="-1" resultid="6791" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1158" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7903" />
                    <RANKING order="2" place="2" resultid="7608" />
                    <RANKING order="3" place="3" resultid="8309" />
                    <RANKING order="4" place="4" resultid="8001" />
                    <RANKING order="5" place="5" resultid="9324" />
                    <RANKING order="6" place="6" resultid="7461" />
                    <RANKING order="7" place="7" resultid="8015" />
                    <RANKING order="8" place="8" resultid="8029" />
                    <RANKING order="9" place="9" resultid="7974" />
                    <RANKING order="10" place="10" resultid="8022" />
                    <RANKING order="11" place="11" resultid="6965" />
                    <RANKING order="12" place="12" resultid="8520" />
                    <RANKING order="13" place="13" resultid="8550" />
                    <RANKING order="14" place="14" resultid="7980" />
                    <RANKING order="15" place="15" resultid="9014" />
                    <RANKING order="16" place="16" resultid="9458" />
                    <RANKING order="17" place="17" resultid="7340" />
                    <RANKING order="18" place="18" resultid="9417" />
                    <RANKING order="19" place="19" resultid="9444" />
                    <RANKING order="20" place="20" resultid="9392" />
                    <RANKING order="21" place="21" resultid="9423" />
                    <RANKING order="22" place="22" resultid="8805" />
                    <RANKING order="23" place="23" resultid="7791" />
                    <RANKING order="24" place="24" resultid="9027" />
                    <RANKING order="25" place="25" resultid="7375" />
                    <RANKING order="26" place="-1" resultid="7915" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1159" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6896" />
                    <RANKING order="2" place="2" resultid="6819" />
                    <RANKING order="3" place="3" resultid="7910" />
                    <RANKING order="4" place="4" resultid="7842" />
                    <RANKING order="5" place="5" resultid="7886" />
                    <RANKING order="6" place="6" resultid="7300" />
                    <RANKING order="7" place="7" resultid="9293" />
                    <RANKING order="8" place="8" resultid="8606" />
                    <RANKING order="9" place="9" resultid="8784" />
                    <RANKING order="10" place="10" resultid="7961" />
                    <RANKING order="11" place="11" resultid="8465" />
                    <RANKING order="12" place="12" resultid="9439" />
                    <RANKING order="13" place="13" resultid="8773" />
                    <RANKING order="14" place="14" resultid="8492" />
                    <RANKING order="15" place="15" resultid="7956" />
                    <RANKING order="16" place="16" resultid="9451" />
                    <RANKING order="17" place="17" resultid="8477" />
                    <RANKING order="18" place="18" resultid="6978" />
                    <RANKING order="19" place="19" resultid="8496" />
                    <RANKING order="20" place="20" resultid="7184" />
                    <RANKING order="21" place="21" resultid="8823" />
                    <RANKING order="22" place="-1" resultid="7848" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1160" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8339" />
                    <RANKING order="2" place="2" resultid="9111" />
                    <RANKING order="3" place="3" resultid="7412" />
                    <RANKING order="4" place="4" resultid="6908" />
                    <RANKING order="5" place="5" resultid="9091" />
                    <RANKING order="6" place="6" resultid="9398" />
                    <RANKING order="7" place="7" resultid="9098" />
                    <RANKING order="8" place="8" resultid="7345" />
                    <RANKING order="9" place="9" resultid="7058" />
                    <RANKING order="10" place="10" resultid="7385" />
                    <RANKING order="11" place="11" resultid="7389" />
                    <RANKING order="12" place="12" resultid="9055" />
                    <RANKING order="13" place="-1" resultid="7837" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1161" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7890" />
                    <RANKING order="2" place="2" resultid="7894" />
                    <RANKING order="3" place="3" resultid="8921" />
                    <RANKING order="4" place="4" resultid="7294" />
                    <RANKING order="5" place="5" resultid="8380" />
                    <RANKING order="6" place="6" resultid="8673" />
                    <RANKING order="7" place="7" resultid="8942" />
                    <RANKING order="8" place="8" resultid="9315" />
                    <RANKING order="9" place="9" resultid="8777" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1162" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8363" />
                    <RANKING order="2" place="2" resultid="7206" />
                    <RANKING order="3" place="3" resultid="9521" />
                    <RANKING order="4" place="4" resultid="9545" />
                    <RANKING order="5" place="5" resultid="9188" />
                    <RANKING order="6" place="6" resultid="9497" />
                    <RANKING order="7" place="7" resultid="9582" />
                    <RANKING order="8" place="8" resultid="9537" />
                    <RANKING order="9" place="9" resultid="9551" />
                    <RANKING order="10" place="10" resultid="7562" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10535" daytime="17:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10536" daytime="17:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10537" daytime="17:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10538" daytime="17:42" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10539" daytime="17:46" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10540" daytime="17:48" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10541" daytime="17:50" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10542" daytime="17:52" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10543" daytime="17:54" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10544" daytime="17:56" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="10545" daytime="17:58" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="10546" daytime="18:00" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="10547" daytime="18:04" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="10548" daytime="18:06" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="10549" daytime="18:08" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="10550" daytime="18:10" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="10551" daytime="18:12" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="10552" daytime="18:12" number="18" order="18" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1163" daytime="18:16" gender="F" number="15" order="5" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1164" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8272" />
                    <RANKING order="2" place="2" resultid="8591" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1165" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7692" />
                    <RANKING order="2" place="2" resultid="7762" />
                    <RANKING order="3" place="3" resultid="8514" />
                    <RANKING order="4" place="4" resultid="7105" />
                    <RANKING order="5" place="-1" resultid="8647" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1166" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9182" />
                    <RANKING order="2" place="2" resultid="8986" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1167" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7867" />
                    <RANKING order="2" place="2" resultid="8556" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1168" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8901" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1169" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7566" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1170" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10553" daytime="18:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10554" daytime="18:20" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1171" daytime="18:26" gender="M" number="16" order="6" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1172" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7508" />
                    <RANKING order="2" place="2" resultid="8217" />
                    <RANKING order="3" place="3" resultid="7720" />
                    <RANKING order="4" place="4" resultid="8620" />
                    <RANKING order="5" place="-1" resultid="8124" />
                    <RANKING order="6" place="-1" resultid="9192" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1173" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7629" />
                    <RANKING order="2" place="2" resultid="9140" />
                    <RANKING order="3" place="3" resultid="9274" />
                    <RANKING order="4" place="4" resultid="7664" />
                    <RANKING order="5" place="5" resultid="7468" />
                    <RANKING order="6" place="6" resultid="9199" />
                    <RANKING order="7" place="7" resultid="8043" />
                    <RANKING order="8" place="8" resultid="8633" />
                    <RANKING order="9" place="9" resultid="8564" />
                    <RANKING order="10" place="10" resultid="8294" />
                    <RANKING order="11" place="-1" resultid="8993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1174" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7482" />
                    <RANKING order="2" place="2" resultid="7776" />
                    <RANKING order="3" place="3" resultid="9147" />
                    <RANKING order="4" place="4" resultid="7615" />
                    <RANKING order="5" place="5" resultid="9013" />
                    <RANKING order="6" place="-1" resultid="7288" />
                    <RANKING order="7" place="-1" resultid="9248" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1175" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7587" />
                    <RANKING order="2" place="2" resultid="7672" />
                    <RANKING order="3" place="3" resultid="8346" />
                    <RANKING order="4" place="4" resultid="6954" />
                    <RANKING order="5" place="5" resultid="7305" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1176" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7713" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1177" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7426" />
                    <RANKING order="2" place="2" resultid="6936" />
                    <RANKING order="3" place="3" resultid="8892" />
                    <RANKING order="4" place="4" resultid="7440" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1178" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8407" />
                    <RANKING order="2" place="2" resultid="7420" />
                    <RANKING order="3" place="3" resultid="9570" />
                    <RANKING order="4" place="4" resultid="9383" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10555" daytime="18:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10556" daytime="18:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10557" daytime="18:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10558" daytime="18:38" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1179" daytime="18:42" gender="F" number="17" order="7" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1180" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8571" />
                    <RANKING order="2" place="2" resultid="9267" />
                    <RANKING order="3" place="3" resultid="9212" />
                    <RANKING order="4" place="4" resultid="8654" />
                    <RANKING order="5" place="5" resultid="7047" />
                    <RANKING order="6" place="6" resultid="7734" />
                    <RANKING order="7" place="7" resultid="7158" />
                    <RANKING order="8" place="8" resultid="9410" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1181" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8332" />
                    <RANKING order="2" place="2" resultid="8071" />
                    <RANKING order="3" place="3" resultid="9133" />
                    <RANKING order="4" place="4" resultid="8597" />
                    <RANKING order="5" place="5" resultid="7488" />
                    <RANKING order="6" place="6" resultid="8717" />
                    <RANKING order="7" place="7" resultid="7123" />
                    <RANKING order="8" place="8" resultid="8402" />
                    <RANKING order="9" place="9" resultid="9356" />
                    <RANKING order="10" place="10" resultid="6586" />
                    <RANKING order="11" place="-1" resultid="9403" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1182" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8872" />
                    <RANKING order="2" place="2" resultid="8300" />
                    <RANKING order="3" place="3" resultid="9219" />
                    <RANKING order="4" place="4" resultid="7924" />
                    <RANKING order="5" place="5" resultid="9234" />
                    <RANKING order="6" place="6" resultid="8693" />
                    <RANKING order="7" place="7" resultid="6995" />
                    <RANKING order="8" place="8" resultid="6859" />
                    <RANKING order="9" place="9" resultid="8535" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1183" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7311" />
                    <RANKING order="2" place="2" resultid="7880" />
                    <RANKING order="3" place="3" resultid="7941" />
                    <RANKING order="4" place="4" resultid="7936" />
                    <RANKING order="5" place="5" resultid="6838" />
                    <RANKING order="6" place="6" resultid="7447" />
                    <RANKING order="7" place="7" resultid="7523" />
                    <RANKING order="8" place="8" resultid="7317" />
                    <RANKING order="9" place="-1" resultid="9065" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1184" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8251" />
                    <RANKING order="2" place="2" resultid="7643" />
                    <RANKING order="3" place="3" resultid="8997" />
                    <RANKING order="4" place="4" resultid="9105" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1185" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7179" />
                    <RANKING order="2" place="2" resultid="9364" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8458" />
                    <RANKING order="2" place="2" resultid="9532" />
                    <RANKING order="3" place="3" resultid="7581" />
                    <RANKING order="4" place="4" resultid="8896" />
                    <RANKING order="5" place="5" resultid="9525" />
                    <RANKING order="6" place="6" resultid="8879" />
                    <RANKING order="7" place="7" resultid="9502" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10560" daytime="18:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10561" daytime="18:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10562" daytime="18:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10563" daytime="18:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10564" daytime="18:48" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10565" daytime="18:50" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1187" daytime="18:52" gender="M" number="18" order="8" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1188" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7018" />
                    <RANKING order="2" place="2" resultid="6932" />
                    <RANKING order="3" place="3" resultid="7252" />
                    <RANKING order="4" place="4" resultid="8619" />
                    <RANKING order="5" place="5" resultid="7116" />
                    <RANKING order="6" place="6" resultid="7755" />
                    <RANKING order="7" place="7" resultid="8794" />
                    <RANKING order="8" place="8" resultid="8230" />
                    <RANKING order="9" place="9" resultid="8660" />
                    <RANKING order="10" place="10" resultid="9434" />
                    <RANKING order="11" place="11" resultid="9330" />
                    <RANKING order="12" place="12" resultid="8723" />
                    <RANKING order="13" place="13" resultid="7379" />
                    <RANKING order="14" place="14" resultid="8813" />
                    <RANKING order="15" place="15" resultid="7502" />
                    <RANKING order="16" place="16" resultid="8818" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1189" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6852" />
                    <RANKING order="2" place="2" resultid="6983" />
                    <RANKING order="3" place="3" resultid="8092" />
                    <RANKING order="4" place="4" resultid="9162" />
                    <RANKING order="5" place="5" resultid="9006" />
                    <RANKING order="6" place="6" resultid="7454" />
                    <RANKING order="7" place="7" resultid="6927" />
                    <RANKING order="8" place="8" resultid="8501" />
                    <RANKING order="9" place="9" resultid="6580" />
                    <RANKING order="10" place="10" resultid="7685" />
                    <RANKING order="11" place="11" resultid="9168" />
                    <RANKING order="12" place="12" resultid="7225" />
                    <RANKING order="13" place="13" resultid="8701" />
                    <RANKING order="14" place="14" resultid="9350" />
                    <RANKING order="15" place="15" resultid="7783" />
                    <RANKING order="16" place="16" resultid="8686" />
                    <RANKING order="17" place="17" resultid="8577" />
                    <RANKING order="18" place="18" resultid="9376" />
                    <RANKING order="19" place="19" resultid="7165" />
                    <RANKING order="20" place="20" resultid="7245" />
                    <RANKING order="21" place="21" resultid="8706" />
                    <RANKING order="22" place="22" resultid="7474" />
                    <RANKING order="23" place="23" resultid="8563" />
                    <RANKING order="24" place="24" resultid="8767" />
                    <RANKING order="25" place="25" resultid="6885" />
                    <RANKING order="26" place="26" resultid="9070" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1190" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8549" />
                    <RANKING order="2" place="2" resultid="9176" />
                    <RANKING order="3" place="3" resultid="9336" />
                    <RANKING order="4" place="4" resultid="8936" />
                    <RANKING order="5" place="5" resultid="7368" />
                    <RANKING order="6" place="6" resultid="7973" />
                    <RANKING order="7" place="7" resultid="9457" />
                    <RANKING order="8" place="8" resultid="7374" />
                    <RANKING order="9" place="9" resultid="9391" />
                    <RANKING order="10" place="10" resultid="7339" />
                    <RANKING order="11" place="11" resultid="8519" />
                    <RANKING order="12" place="12" resultid="8804" />
                    <RANKING order="13" place="13" resultid="9026" />
                    <RANKING order="14" place="-1" resultid="7790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1191" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8914" />
                    <RANKING order="2" place="2" resultid="8375" />
                    <RANKING order="3" place="3" resultid="8395" />
                    <RANKING order="4" place="4" resultid="7946" />
                    <RANKING order="5" place="5" resultid="8783" />
                    <RANKING order="6" place="6" resultid="6915" />
                    <RANKING order="7" place="7" resultid="8464" />
                    <RANKING order="8" place="8" resultid="8476" />
                    <RANKING order="9" place="9" resultid="9450" />
                    <RANKING order="10" place="10" resultid="6977" />
                    <RANKING order="11" place="11" resultid="7183" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1192" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6947" />
                    <RANKING order="2" place="2" resultid="7852" />
                    <RANKING order="3" place="3" resultid="8338" />
                    <RANKING order="4" place="4" resultid="8960" />
                    <RANKING order="5" place="5" resultid="7057" />
                    <RANKING order="6" place="6" resultid="6989" />
                    <RANKING order="7" place="7" resultid="9097" />
                    <RANKING order="8" place="8" resultid="8505" />
                    <RANKING order="9" place="9" resultid="9054" />
                    <RANKING order="10" place="-1" resultid="6921" />
                    <RANKING order="11" place="-1" resultid="8291" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1193" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7899" />
                    <RANKING order="2" place="2" resultid="6560" />
                    <RANKING order="3" place="3" resultid="7622" />
                    <RANKING order="4" place="4" resultid="7531" />
                    <RANKING order="5" place="-1" resultid="8391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1194" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9513" />
                    <RANKING order="2" place="2" resultid="6824" />
                    <RANKING order="3" place="3" resultid="9520" />
                    <RANKING order="4" place="4" resultid="7201" />
                    <RANKING order="5" place="5" resultid="9600" />
                    <RANKING order="6" place="6" resultid="9507" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10566" daytime="18:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10567" daytime="18:54" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10568" daytime="18:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10569" daytime="18:58" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10570" daytime="19:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10571" daytime="19:02" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10572" daytime="19:04" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10573" daytime="19:06" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10574" daytime="19:08" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10575" daytime="19:08" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1195" daytime="19:20" gender="F" number="19" order="10" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1196" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8410" />
                    <RANKING order="2" place="2" resultid="9463" />
                    <RANKING order="3" place="3" resultid="7802" />
                    <RANKING order="4" place="4" resultid="8745" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10576" daytime="19:20" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1197" daytime="19:32" gender="F" number="20" order="11" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1198" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8409" />
                    <RANKING order="2" place="2" resultid="7801" />
                    <RANKING order="3" place="3" resultid="9462" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10577" daytime="19:32" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1199" daytime="19:44" gender="F" number="21" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1200" agemax="19" agemin="17" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1201" daytime="19:44" gender="F" number="22" order="13" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1202" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9609" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10578" daytime="19:44" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1203" daytime="19:54" gender="M" number="23" order="14" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1204" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8421" />
                    <RANKING order="2" place="2" resultid="7809" />
                    <RANKING order="3" place="3" resultid="9472" />
                    <RANKING order="4" place="4" resultid="7515" />
                    <RANKING order="5" place="5" resultid="8749" />
                    <RANKING order="6" place="6" resultid="7257" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10579" daytime="19:54" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1205" daytime="20:06" gender="M" number="24" order="15" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1206" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8419" />
                    <RANKING order="2" place="2" resultid="7807" />
                    <RANKING order="3" place="3" resultid="9470" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10580" daytime="20:06" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1207" daytime="20:18" gender="M" number="25" order="16" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1208" agemax="19" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8420" />
                    <RANKING order="2" place="2" resultid="7808" />
                    <RANKING order="3" place="3" resultid="7514" />
                    <RANKING order="4" place="4" resultid="9471" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10581" daytime="20:18" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1209" daytime="20:28" gender="M" number="26" order="17" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1210" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9612" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10582" daytime="20:28" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2025-04-12" daytime="08:55" endtime="13:27" number="3" officialmeeting="08:00" status="OFFICIAL" warmupfrom="07:30" warmupuntil="08:30">
          <EVENTS>
            <EVENT eventid="1211" daytime="08:56" gender="F" number="27" order="1" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1212" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8193" />
                    <RANKING order="2" place="2" resultid="8574" />
                    <RANKING order="3" place="3" resultid="8146" />
                    <RANKING order="4" place="4" resultid="9268" />
                    <RANKING order="5" place="5" resultid="8226" />
                    <RANKING order="6" place="6" resultid="8357" />
                    <RANKING order="7" place="7" resultid="8656" />
                    <RANKING order="8" place="8" resultid="7048" />
                    <RANKING order="9" place="9" resultid="7736" />
                    <RANKING order="10" place="10" resultid="9049" />
                    <RANKING order="11" place="11" resultid="8317" />
                    <RANKING order="12" place="12" resultid="9215" />
                    <RANKING order="13" place="13" resultid="9243" />
                    <RANKING order="14" place="14" resultid="9431" />
                    <RANKING order="15" place="15" resultid="9413" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1213" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8067" />
                    <RANKING order="2" place="2" resultid="8074" />
                    <RANKING order="3" place="3" resultid="8335" />
                    <RANKING order="4" place="4" resultid="7694" />
                    <RANKING order="5" place="5" resultid="8246" />
                    <RANKING order="6" place="6" resultid="8081" />
                    <RANKING order="7" place="7" resultid="9136" />
                    <RANKING order="8" place="8" resultid="8515" />
                    <RANKING order="9" place="9" resultid="7764" />
                    <RANKING order="10" place="10" resultid="8405" />
                    <RANKING order="11" place="11" resultid="9034" />
                    <RANKING order="12" place="12" resultid="9359" />
                    <RANKING order="13" place="13" resultid="9406" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1214" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8875" />
                    <RANKING order="2" place="2" resultid="7701" />
                    <RANKING order="3" place="3" resultid="8303" />
                    <RANKING order="4" place="4" resultid="7875" />
                    <RANKING order="5" place="5" resultid="9220" />
                    <RANKING order="6" place="6" resultid="9235" />
                    <RANKING order="7" place="7" resultid="8695" />
                    <RANKING order="8" place="8" resultid="6869" />
                    <RANKING order="9" place="9" resultid="8537" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1215" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7937" />
                    <RANKING order="2" place="2" resultid="7881" />
                    <RANKING order="3" place="3" resultid="7312" />
                    <RANKING order="4" place="4" resultid="7823" />
                    <RANKING order="5" place="5" resultid="7602" />
                    <RANKING order="6" place="6" resultid="6839" />
                    <RANKING order="7" place="7" resultid="7526" />
                    <RANKING order="8" place="-1" resultid="7942" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1216" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8253" />
                    <RANKING order="2" place="2" resultid="7645" />
                    <RANKING order="3" place="3" resultid="7096" />
                    <RANKING order="4" place="4" resultid="9000" />
                    <RANKING order="5" place="5" resultid="9107" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1217" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7856" />
                    <RANKING order="2" place="2" resultid="7180" />
                    <RANKING order="3" place="3" resultid="9365" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1218" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8459" />
                    <RANKING order="2" place="2" resultid="9533" />
                    <RANKING order="3" place="3" resultid="7582" />
                    <RANKING order="4" place="4" resultid="8897" />
                    <RANKING order="5" place="5" resultid="9528" />
                    <RANKING order="6" place="6" resultid="8880" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10583" daytime="08:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10584" daytime="08:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10585" daytime="09:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10586" daytime="09:04" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10587" daytime="09:06" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10588" daytime="09:08" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10589" daytime="09:10" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1219" daytime="09:14" gender="M" number="28" order="2" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1220" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8287" />
                    <RANKING order="2" place="2" resultid="8179" />
                    <RANKING order="3" place="3" resultid="8212" />
                    <RANKING order="4" place="4" resultid="9195" />
                    <RANKING order="5" place="5" resultid="7756" />
                    <RANKING order="6" place="6" resultid="8621" />
                    <RANKING order="7" place="7" resultid="6933" />
                    <RANKING order="8" place="8" resultid="7119" />
                    <RANKING order="9" place="9" resultid="8232" />
                    <RANKING order="10" place="10" resultid="8173" />
                    <RANKING order="11" place="11" resultid="8726" />
                    <RANKING order="12" place="12" resultid="8816" />
                    <RANKING order="13" place="13" resultid="9255" />
                    <RANKING order="14" place="14" resultid="7382" />
                    <RANKING order="15" place="-1" resultid="9332" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1221" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7750" />
                    <RANKING order="2" place="2" resultid="8095" />
                    <RANKING order="3" place="3" resultid="6855" />
                    <RANKING order="4" place="4" resultid="6984" />
                    <RANKING order="5" place="5" resultid="9164" />
                    <RANKING order="6" place="6" resultid="8052" />
                    <RANKING order="7" place="7" resultid="6928" />
                    <RANKING order="8" place="8" resultid="7652" />
                    <RANKING order="9" place="9" resultid="8281" />
                    <RANKING order="10" place="10" resultid="9008" />
                    <RANKING order="11" place="11" resultid="7686" />
                    <RANKING order="12" place="12" resultid="8114" />
                    <RANKING order="13" place="13" resultid="9171" />
                    <RANKING order="14" place="14" resultid="6582" />
                    <RANKING order="15" place="15" resultid="7226" />
                    <RANKING order="16" place="16" resultid="8635" />
                    <RANKING order="17" place="17" resultid="9352" />
                    <RANKING order="18" place="18" resultid="6736" />
                    <RANKING order="19" place="19" resultid="7786" />
                    <RANKING order="20" place="20" resultid="8580" />
                    <RANKING order="21" place="21" resultid="9043" />
                    <RANKING order="22" place="22" resultid="7248" />
                    <RANKING order="23" place="23" resultid="7477" />
                    <RANKING order="24" place="24" resultid="6888" />
                    <RANKING order="25" place="-1" resultid="6779" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1222" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8552" />
                    <RANKING order="2" place="2" resultid="9177" />
                    <RANKING order="3" place="3" resultid="8938" />
                    <RANKING order="4" place="4" resultid="8017" />
                    <RANKING order="5" place="5" resultid="9337" />
                    <RANKING order="6" place="6" resultid="7369" />
                    <RANKING order="7" place="7" resultid="7976" />
                    <RANKING order="8" place="8" resultid="8948" />
                    <RANKING order="9" place="9" resultid="7377" />
                    <RANKING order="10" place="10" resultid="9394" />
                    <RANKING order="11" place="11" resultid="7793" />
                    <RANKING order="12" place="-1" resultid="7982" />
                    <RANKING order="13" place="-1" resultid="8522" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1223" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8915" />
                    <RANKING order="2" place="2" resultid="8376" />
                    <RANKING order="3" place="3" resultid="8396" />
                    <RANKING order="4" place="4" resultid="7301" />
                    <RANKING order="5" place="5" resultid="6917" />
                    <RANKING order="6" place="6" resultid="7947" />
                    <RANKING order="7" place="7" resultid="8786" />
                    <RANKING order="8" place="8" resultid="6979" />
                    <RANKING order="9" place="-1" resultid="7843" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1224" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8268" />
                    <RANKING order="2" place="2" resultid="7854" />
                    <RANKING order="3" place="3" resultid="6949" />
                    <RANKING order="4" place="4" resultid="7435" />
                    <RANKING order="5" place="5" resultid="8961" />
                    <RANKING order="6" place="6" resultid="7680" />
                    <RANKING order="7" place="7" resultid="8507" />
                    <RANKING order="8" place="8" resultid="9056" />
                    <RANKING order="9" place="-1" resultid="7060" />
                    <RANKING order="10" place="-1" resultid="6922" />
                    <RANKING order="11" place="-1" resultid="8341" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1225" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7900" />
                    <RANKING order="2" place="2" resultid="6561" />
                    <RANKING order="3" place="3" resultid="7624" />
                    <RANKING order="4" place="4" resultid="7532" />
                    <RANKING order="5" place="-1" resultid="8392" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1226" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7970" />
                    <RANKING order="2" place="2" resultid="9515" />
                    <RANKING order="3" place="3" resultid="6825" />
                    <RANKING order="4" place="4" resultid="9566" />
                    <RANKING order="5" place="5" resultid="9538" />
                    <RANKING order="6" place="6" resultid="9601" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10590" daytime="09:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10591" daytime="09:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10592" daytime="09:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10593" daytime="09:22" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10594" daytime="09:24" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10595" daytime="09:28" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10596" daytime="09:30" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10597" daytime="09:32" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10598" daytime="09:34" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10599" daytime="09:36" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1227" daytime="09:40" gender="F" number="29" order="3" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1228" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8263" />
                    <RANKING order="2" place="2" resultid="8273" />
                    <RANKING order="3" place="3" resultid="8573" />
                    <RANKING order="4" place="4" resultid="9242" />
                    <RANKING order="5" place="5" resultid="8356" />
                    <RANKING order="6" place="6" resultid="8593" />
                    <RANKING order="7" place="7" resultid="8738" />
                    <RANKING order="8" place="8" resultid="8206" />
                    <RANKING order="9" place="9" resultid="7134" />
                    <RANKING order="10" place="10" resultid="8192" />
                    <RANKING order="11" place="11" resultid="9214" />
                    <RANKING order="12" place="12" resultid="9605" />
                    <RANKING order="13" place="13" resultid="8655" />
                    <RANKING order="14" place="14" resultid="8790" />
                    <RANKING order="15" place="15" resultid="7160" />
                    <RANKING order="16" place="16" resultid="8526" />
                    <RANKING order="17" place="17" resultid="7363" />
                    <RANKING order="18" place="18" resultid="9412" />
                    <RANKING order="19" place="19" resultid="8667" />
                    <RANKING order="20" place="-1" resultid="9430" />
                    <RANKING order="21" place="-1" resultid="8257" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1229" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6880" />
                    <RANKING order="2" place="2" resultid="8599" />
                    <RANKING order="3" place="3" resultid="8086" />
                    <RANKING order="4" place="4" resultid="8326" />
                    <RANKING order="5" place="5" resultid="8080" />
                    <RANKING order="6" place="6" resultid="8487" />
                    <RANKING order="7" place="7" resultid="6874" />
                    <RANKING order="8" place="8" resultid="9371" />
                    <RANKING order="9" place="9" resultid="8245" />
                    <RANKING order="10" place="10" resultid="8334" />
                    <RANKING order="11" place="11" resultid="7537" />
                    <RANKING order="12" place="12" resultid="7007" />
                    <RANKING order="13" place="13" resultid="7490" />
                    <RANKING order="14" place="14" resultid="9135" />
                    <RANKING order="15" place="15" resultid="7013" />
                    <RANKING order="16" place="16" resultid="9283" />
                    <RANKING order="17" place="17" resultid="8404" />
                    <RANKING order="18" place="18" resultid="6588" />
                    <RANKING order="19" place="19" resultid="9289" />
                    <RANKING order="20" place="20" resultid="7106" />
                    <RANKING order="21" place="21" resultid="9405" />
                    <RANKING order="22" place="22" resultid="8719" />
                    <RANKING order="23" place="23" resultid="9358" />
                    <RANKING order="24" place="-1" resultid="6701" />
                    <RANKING order="25" place="-1" resultid="9155" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1230" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6574" />
                    <RANKING order="2" place="2" resultid="6567" />
                    <RANKING order="3" place="3" resultid="7100" />
                    <RANKING order="4" place="4" resultid="7926" />
                    <RANKING order="5" place="5" resultid="7989" />
                    <RANKING order="6" place="6" resultid="7196" />
                    <RANKING order="7" place="7" resultid="7001" />
                    <RANKING order="8" place="8" resultid="7994" />
                    <RANKING order="9" place="9" resultid="9301" />
                    <RANKING order="10" place="10" resultid="9588" />
                    <RANKING order="11" place="11" resultid="7596" />
                    <RANKING order="12" place="12" resultid="8614" />
                    <RANKING order="13" place="13" resultid="7082" />
                    <RANKING order="14" place="14" resultid="7220" />
                    <RANKING order="15" place="15" resultid="6863" />
                    <RANKING order="16" place="16" resultid="9309" />
                    <RANKING order="17" place="17" resultid="8800" />
                    <RANKING order="18" place="18" resultid="6868" />
                    <RANKING order="19" place="19" resultid="8536" />
                    <RANKING order="20" place="20" resultid="7557" />
                    <RANKING order="21" place="-1" resultid="8302" />
                    <RANKING order="22" place="-1" resultid="7153" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1231" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7829" />
                    <RANKING order="2" place="2" resultid="6829" />
                    <RANKING order="3" place="3" resultid="7868" />
                    <RANKING order="4" place="4" resultid="7952" />
                    <RANKING order="5" place="5" resultid="7319" />
                    <RANKING order="6" place="6" resultid="7216" />
                    <RANKING order="7" place="7" resultid="8557" />
                    <RANKING order="8" place="8" resultid="7449" />
                    <RANKING order="9" place="9" resultid="6943" />
                    <RANKING order="10" place="10" resultid="7525" />
                    <RANKING order="11" place="11" resultid="9066" />
                    <RANKING order="12" place="-1" resultid="6646" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1232" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8999" />
                    <RANKING order="2" place="2" resultid="7089" />
                    <RANKING order="3" place="3" resultid="8252" />
                    <RANKING order="4" place="4" resultid="7095" />
                    <RANKING order="5" place="5" resultid="7352" />
                    <RANKING order="6" place="6" resultid="6961" />
                    <RANKING order="7" place="7" resultid="7129" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1233" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6833" />
                    <RANKING order="2" place="2" resultid="9085" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1234" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7405" />
                    <RANKING order="2" place="2" resultid="9527" />
                    <RANKING order="3" place="3" resultid="9578" />
                    <RANKING order="4" place="4" resultid="9504" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10600" daytime="09:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10601" daytime="09:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10602" daytime="09:42" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10603" daytime="09:44" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10604" daytime="09:46" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10605" daytime="09:48" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10606" daytime="09:50" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10607" daytime="09:50" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10608" daytime="09:52" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10609" daytime="09:54" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1235" daytime="09:56" gender="M" number="30" order="4" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1236" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7510" />
                    <RANKING order="2" place="2" resultid="8387" />
                    <RANKING order="3" place="3" resultid="7030" />
                    <RANKING order="4" place="4" resultid="7148" />
                    <RANKING order="5" place="5" resultid="9194" />
                    <RANKING order="6" place="6" resultid="8166" />
                    <RANKING order="7" place="7" resultid="7358" />
                    <RANKING order="8" place="8" resultid="8662" />
                    <RANKING order="9" place="9" resultid="8132" />
                    <RANKING order="10" place="10" resultid="7173" />
                    <RANKING order="11" place="11" resultid="8585" />
                    <RANKING order="12" place="12" resultid="7020" />
                    <RANKING order="13" place="13" resultid="8186" />
                    <RANKING order="14" place="14" resultid="7324" />
                    <RANKING order="15" place="15" resultid="9343" />
                    <RANKING order="16" place="16" resultid="7112" />
                    <RANKING order="17" place="17" resultid="8159" />
                    <RANKING order="18" place="18" resultid="8954" />
                    <RANKING order="19" place="19" resultid="8138" />
                    <RANKING order="20" place="20" resultid="8482" />
                    <RANKING order="21" place="21" resultid="8744" />
                    <RANKING order="22" place="22" resultid="7042" />
                    <RANKING order="23" place="23" resultid="7504" />
                    <RANKING order="24" place="23" resultid="8725" />
                    <RANKING order="25" place="25" resultid="9261" />
                    <RANKING order="26" place="26" resultid="7053" />
                    <RANKING order="27" place="27" resultid="7381" />
                    <RANKING order="28" place="28" resultid="7118" />
                    <RANKING order="29" place="29" resultid="7254" />
                    <RANKING order="30" place="30" resultid="9254" />
                    <RANKING order="31" place="31" resultid="8172" />
                    <RANKING order="32" place="32" resultid="9436" />
                    <RANKING order="33" place="33" resultid="8763" />
                    <RANKING order="34" place="34" resultid="8815" />
                    <RANKING order="35" place="35" resultid="8820" />
                    <RANKING order="36" place="-1" resultid="8125" />
                    <RANKING order="37" place="-1" resultid="8218" />
                    <RANKING order="38" place="-1" resultid="8731" />
                    <RANKING order="39" place="-1" resultid="6743" />
                    <RANKING order="40" place="-1" resultid="9227" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1237" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6903" />
                    <RANKING order="2" place="2" resultid="8239" />
                    <RANKING order="3" place="3" resultid="8626" />
                    <RANKING order="4" place="4" resultid="7142" />
                    <RANKING order="5" place="5" resultid="8094" />
                    <RANKING order="6" place="6" resultid="7456" />
                    <RANKING order="7" place="7" resultid="8038" />
                    <RANKING order="8" place="8" resultid="6854" />
                    <RANKING order="9" place="9" resultid="8051" />
                    <RANKING order="10" place="10" resultid="9275" />
                    <RANKING order="11" place="11" resultid="8641" />
                    <RANKING order="12" place="12" resultid="7231" />
                    <RANKING order="13" place="12" resultid="7543" />
                    <RANKING order="14" place="14" resultid="8369" />
                    <RANKING order="15" place="15" resultid="7469" />
                    <RANKING order="16" place="16" resultid="8472" />
                    <RANKING order="17" place="17" resultid="7063" />
                    <RANKING order="18" place="18" resultid="9207" />
                    <RANKING order="19" place="19" resultid="9170" />
                    <RANKING order="20" place="20" resultid="8687" />
                    <RANKING order="21" place="21" resultid="9163" />
                    <RANKING order="22" place="22" resultid="7240" />
                    <RANKING order="23" place="23" resultid="7167" />
                    <RANKING order="24" place="24" resultid="8502" />
                    <RANKING order="25" place="25" resultid="7549" />
                    <RANKING order="26" place="26" resultid="7247" />
                    <RANKING order="27" place="26" resultid="8296" />
                    <RANKING order="28" place="28" resultid="8101" />
                    <RANKING order="29" place="29" resultid="7329" />
                    <RANKING order="30" place="30" resultid="8565" />
                    <RANKING order="31" place="31" resultid="6973" />
                    <RANKING order="32" place="32" resultid="8634" />
                    <RANKING order="33" place="33" resultid="8702" />
                    <RANKING order="34" place="34" resultid="9378" />
                    <RANKING order="35" place="35" resultid="7236" />
                    <RANKING order="36" place="36" resultid="7476" />
                    <RANKING order="37" place="37" resultid="6887" />
                    <RANKING order="38" place="38" resultid="7785" />
                    <RANKING order="39" place="39" resultid="9042" />
                    <RANKING order="40" place="40" resultid="8579" />
                    <RANKING order="41" place="41" resultid="8994" />
                    <RANKING order="42" place="42" resultid="9072" />
                    <RANKING order="43" place="43" resultid="8810" />
                    <RANKING order="44" place="44" resultid="8708" />
                    <RANKING order="45" place="45" resultid="8769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1238" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7904" />
                    <RANKING order="2" place="2" resultid="7462" />
                    <RANKING order="3" place="3" resultid="8310" />
                    <RANKING order="4" place="4" resultid="8002" />
                    <RANKING order="5" place="5" resultid="8016" />
                    <RANKING order="6" place="6" resultid="9325" />
                    <RANKING order="7" place="7" resultid="7975" />
                    <RANKING order="8" place="8" resultid="9148" />
                    <RANKING order="9" place="9" resultid="8023" />
                    <RANKING order="10" place="9" resultid="8031" />
                    <RANKING order="11" place="11" resultid="8531" />
                    <RANKING order="12" place="12" resultid="7483" />
                    <RANKING order="13" place="13" resultid="6966" />
                    <RANKING order="14" place="14" resultid="8521" />
                    <RANKING order="15" place="15" resultid="8551" />
                    <RANKING order="16" place="16" resultid="9459" />
                    <RANKING order="17" place="17" resultid="7341" />
                    <RANKING order="18" place="18" resultid="9418" />
                    <RANKING order="19" place="19" resultid="8806" />
                    <RANKING order="20" place="20" resultid="9028" />
                    <RANKING order="21" place="21" resultid="9445" />
                    <RANKING order="22" place="22" resultid="7792" />
                    <RANKING order="23" place="23" resultid="9393" />
                    <RANKING order="24" place="24" resultid="9424" />
                    <RANKING order="25" place="25" resultid="7376" />
                    <RANKING order="26" place="-1" resultid="7917" />
                    <RANKING order="27" place="-1" resultid="7981" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1239" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6897" />
                    <RANKING order="2" place="2" resultid="6820" />
                    <RANKING order="3" place="3" resultid="8347" />
                    <RANKING order="4" place="4" resultid="8785" />
                    <RANKING order="5" place="5" resultid="6955" />
                    <RANKING order="6" place="6" resultid="8774" />
                    <RANKING order="7" place="7" resultid="9294" />
                    <RANKING order="8" place="8" resultid="7306" />
                    <RANKING order="9" place="9" resultid="9440" />
                    <RANKING order="10" place="10" resultid="8466" />
                    <RANKING order="11" place="11" resultid="9452" />
                    <RANKING order="12" place="12" resultid="6916" />
                    <RANKING order="13" place="13" resultid="8493" />
                    <RANKING order="14" place="14" resultid="7957" />
                    <RANKING order="15" place="15" resultid="7931" />
                    <RANKING order="16" place="16" resultid="8478" />
                    <RANKING order="17" place="17" resultid="8497" />
                    <RANKING order="18" place="18" resultid="8824" />
                    <RANKING order="19" place="-1" resultid="7849" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1240" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8340" />
                    <RANKING order="2" place="2" resultid="7413" />
                    <RANKING order="3" place="3" resultid="9112" />
                    <RANKING order="4" place="4" resultid="9399" />
                    <RANKING order="5" place="5" resultid="7575" />
                    <RANKING order="6" place="6" resultid="6909" />
                    <RANKING order="7" place="7" resultid="7853" />
                    <RANKING order="8" place="8" resultid="6948" />
                    <RANKING order="9" place="9" resultid="9099" />
                    <RANKING order="10" place="10" resultid="9092" />
                    <RANKING order="11" place="11" resultid="7346" />
                    <RANKING order="12" place="12" resultid="7059" />
                    <RANKING order="13" place="13" resultid="7390" />
                    <RANKING order="14" place="14" resultid="6990" />
                    <RANKING order="15" place="15" resultid="7386" />
                    <RANKING order="16" place="16" resultid="8506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1241" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7891" />
                    <RANKING order="2" place="2" resultid="7895" />
                    <RANKING order="3" place="3" resultid="8922" />
                    <RANKING order="4" place="4" resultid="8381" />
                    <RANKING order="5" place="5" resultid="6847" />
                    <RANKING order="6" place="6" resultid="8893" />
                    <RANKING order="7" place="7" resultid="6937" />
                    <RANKING order="8" place="8" resultid="7295" />
                    <RANKING order="9" place="9" resultid="8674" />
                    <RANKING order="10" place="10" resultid="9316" />
                    <RANKING order="11" place="11" resultid="7442" />
                    <RANKING order="12" place="12" resultid="8778" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1242" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8364" />
                    <RANKING order="2" place="2" resultid="7207" />
                    <RANKING order="3" place="3" resultid="7408" />
                    <RANKING order="4" place="4" resultid="8306" />
                    <RANKING order="5" place="5" resultid="9522" />
                    <RANKING order="6" place="6" resultid="9514" />
                    <RANKING order="7" place="7" resultid="9119" />
                    <RANKING order="8" place="8" resultid="9583" />
                    <RANKING order="9" place="9" resultid="9320" />
                    <RANKING order="10" place="10" resultid="9546" />
                    <RANKING order="11" place="11" resultid="9498" />
                    <RANKING order="12" place="12" resultid="7191" />
                    <RANKING order="13" place="13" resultid="9571" />
                    <RANKING order="14" place="14" resultid="9385" />
                    <RANKING order="15" place="15" resultid="9508" />
                    <RANKING order="16" place="16" resultid="9552" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10610" daytime="09:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10611" daytime="09:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10612" daytime="10:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10613" daytime="10:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10614" daytime="10:02" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10615" daytime="10:04" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10616" daytime="10:06" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10617" daytime="10:08" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10618" daytime="10:08" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10619" daytime="10:10" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="10620" daytime="10:12" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="10621" daytime="10:14" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="10622" daytime="10:14" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="10623" daytime="10:16" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="10624" daytime="10:18" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="10625" daytime="10:20" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="10626" daytime="10:20" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="10627" daytime="10:22" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="10628" daytime="10:24" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="10793" daytime="10:24" number="20" order="20" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1243" daytime="10:42" gender="X" number="31" order="6" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1244" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7818" />
                    <RANKING order="2" place="2" resultid="8435" />
                    <RANKING order="3" place="3" resultid="9486" />
                    <RANKING order="4" place="4" resultid="8453" />
                    <RANKING order="5" place="5" resultid="9494" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10629" daytime="10:42" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1245" daytime="10:48" gender="X" number="32" order="7" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1246" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8436" />
                    <RANKING order="2" place="2" resultid="8454" />
                    <RANKING order="3" place="3" resultid="7395" />
                    <RANKING order="4" place="4" resultid="7819" />
                    <RANKING order="5" place="5" resultid="8756" />
                    <RANKING order="6" place="6" resultid="7078" />
                    <RANKING order="7" place="7" resultid="6892" />
                    <RANKING order="8" place="8" resultid="9487" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10630" daytime="10:48" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1247" daytime="10:56" gender="X" number="33" order="8" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1248" agemax="-1" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7817" />
                    <RANKING order="2" place="2" resultid="8434" />
                    <RANKING order="3" place="3" resultid="7520" />
                    <RANKING order="4" place="4" resultid="9485" />
                    <RANKING order="5" place="5" resultid="9615" />
                    <RANKING order="6" place="6" resultid="9618" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10631" daytime="10:56" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1249" daytime="11:02" gender="F" number="34" order="9" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1250" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8152" />
                    <RANKING order="2" place="2" resultid="8199" />
                    <RANKING order="3" place="3" resultid="8225" />
                    <RANKING order="4" place="4" resultid="8145" />
                    <RANKING order="5" place="5" resultid="9048" />
                    <RANKING order="6" place="6" resultid="8592" />
                    <RANKING order="7" place="7" resultid="9020" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1251" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8066" />
                    <RANKING order="2" place="2" resultid="8108" />
                    <RANKING order="3" place="3" resultid="7659" />
                    <RANKING order="4" place="4" resultid="7743" />
                    <RANKING order="5" place="5" resultid="8073" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1252" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7700" />
                    <RANKING order="2" place="2" resultid="7496" />
                    <RANKING order="3" place="3" resultid="8929" />
                    <RANKING order="4" place="4" resultid="8874" />
                    <RANKING order="5" place="5" resultid="7770" />
                    <RANKING order="6" place="6" resultid="8613" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1253" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7862" />
                    <RANKING order="2" place="-1" resultid="6645" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1254" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8966" />
                    <RANKING order="2" place="2" resultid="7211" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1255" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8681" />
                    <RANKING order="2" place="2" resultid="7567" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1256" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9577" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10632" daytime="11:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10633" daytime="11:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10634" daytime="11:26" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1257" daytime="11:40" gender="M" number="35" order="10" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1258" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7721" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1259" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8037" />
                    <RANKING order="2" place="2" resultid="7630" />
                    <RANKING order="3" place="3" resultid="8974" />
                    <RANKING order="4" place="4" resultid="8044" />
                    <RANKING order="5" place="5" resultid="9007" />
                    <RANKING order="6" place="6" resultid="8059" />
                    <RANKING order="7" place="7" resultid="9200" />
                    <RANKING order="8" place="8" resultid="8280" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1260" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8030" />
                    <RANKING order="2" place="2" resultid="7708" />
                    <RANKING order="3" place="3" resultid="8937" />
                    <RANKING order="4" place="4" resultid="9249" />
                    <RANKING order="5" place="5" resultid="8947" />
                    <RANKING order="6" place="6" resultid="7616" />
                    <RANKING order="7" place="-1" resultid="7916" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1261" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8909" />
                    <RANKING order="2" place="2" resultid="7589" />
                    <RANKING order="3" place="3" resultid="7962" />
                    <RANKING order="4" place="4" resultid="8607" />
                    <RANKING order="5" place="5" resultid="6843" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1262" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7714" />
                    <RANKING order="2" place="2" resultid="8510" />
                    <RANKING order="3" place="-1" resultid="7434" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1263" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7441" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1264" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9384" />
                    <RANKING order="2" place="2" resultid="9565" />
                    <RANKING order="3" place="3" resultid="9558" />
                    <RANKING order="4" place="4" resultid="9594" />
                    <RANKING order="5" place="-1" resultid="7563" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10635" daytime="11:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10636" daytime="12:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10637" daytime="12:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10638" daytime="12:44" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2025-04-12" daytime="15:55" endtime="20:11" number="4" officialmeeting="15:00" status="OFFICIAL" warmupfrom="14:30" warmupuntil="15:30">
          <EVENTS>
            <EVENT eventid="1265" daytime="15:56" gender="F" number="36" order="1" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1266" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8274" />
                    <RANKING order="2" place="2" resultid="8200" />
                    <RANKING order="3" place="3" resultid="8227" />
                    <RANKING order="4" place="4" resultid="9244" />
                    <RANKING order="5" place="4" resultid="9269" />
                    <RANKING order="6" place="6" resultid="8194" />
                    <RANKING order="7" place="7" resultid="7737" />
                    <RANKING order="8" place="8" resultid="7049" />
                    <RANKING order="9" place="9" resultid="9021" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1267" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8068" />
                    <RANKING order="2" place="2" resultid="8247" />
                    <RANKING order="3" place="3" resultid="8327" />
                    <RANKING order="4" place="4" resultid="7765" />
                    <RANKING order="5" place="5" resultid="7695" />
                    <RANKING order="6" place="6" resultid="8516" />
                    <RANKING order="7" place="7" resultid="7539" />
                    <RANKING order="8" place="8" resultid="7125" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1268" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7702" />
                    <RANKING order="2" place="2" resultid="7877" />
                    <RANKING order="3" place="3" resultid="7995" />
                    <RANKING order="4" place="4" resultid="9236" />
                    <RANKING order="5" place="5" resultid="8876" />
                    <RANKING order="6" place="6" resultid="9221" />
                    <RANKING order="7" place="7" resultid="7990" />
                    <RANKING order="8" place="8" resultid="8931" />
                    <RANKING order="9" place="9" resultid="8987" />
                    <RANKING order="10" place="10" resultid="8981" />
                    <RANKING order="11" place="-1" resultid="9302" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1269" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7882" />
                    <RANKING order="2" place="2" resultid="8558" />
                    <RANKING order="3" place="3" resultid="7943" />
                    <RANKING order="4" place="4" resultid="7603" />
                    <RANKING order="5" place="5" resultid="7527" />
                    <RANKING order="6" place="-1" resultid="7284" />
                    <RANKING order="7" place="-1" resultid="6647" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1270" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7646" />
                    <RANKING order="2" place="2" resultid="7400" />
                    <RANKING order="3" place="3" resultid="8903" />
                    <RANKING order="4" place="4" resultid="9108" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1271" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7181" />
                    <RANKING order="2" place="2" resultid="8682" />
                    <RANKING order="3" place="3" resultid="9367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1272" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7583" />
                    <RANKING order="2" place="2" resultid="8881" />
                    <RANKING order="3" place="-1" resultid="9534" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10639" daytime="15:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10640" daytime="16:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10641" daytime="16:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10642" daytime="16:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10643" daytime="16:12" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10644" daytime="16:16" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1273" daytime="16:20" gender="M" number="37" order="2" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1274" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7037" />
                    <RANKING order="2" place="2" resultid="8288" />
                    <RANKING order="3" place="3" resultid="8219" />
                    <RANKING order="4" place="4" resultid="8956" />
                    <RANKING order="5" place="5" resultid="8587" />
                    <RANKING order="6" place="6" resultid="8796" />
                    <RANKING order="7" place="7" resultid="7638" />
                    <RANKING order="8" place="8" resultid="7757" />
                    <RANKING order="9" place="9" resultid="8174" />
                    <RANKING order="10" place="-1" resultid="8213" />
                    <RANKING order="11" place="-1" resultid="9345" />
                    <RANKING order="12" place="-1" resultid="6759" />
                    <RANKING order="13" place="-1" resultid="6744" />
                    <RANKING order="14" place="-1" resultid="9228" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1275" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9142" />
                    <RANKING order="2" place="2" resultid="7653" />
                    <RANKING order="3" place="3" resultid="8115" />
                    <RANKING order="4" place="4" resultid="7751" />
                    <RANKING order="5" place="5" resultid="7729" />
                    <RANKING order="6" place="6" resultid="7666" />
                    <RANKING order="7" place="7" resultid="8282" />
                    <RANKING order="8" place="8" resultid="9165" />
                    <RANKING order="9" place="9" resultid="9172" />
                    <RANKING order="10" place="10" resultid="9009" />
                    <RANKING order="11" place="11" resultid="8636" />
                    <RANKING order="12" place="12" resultid="6929" />
                    <RANKING order="13" place="13" resultid="7687" />
                    <RANKING order="14" place="14" resultid="8689" />
                    <RANKING order="15" place="15" resultid="8703" />
                    <RANKING order="16" place="16" resultid="7550" />
                    <RANKING order="17" place="17" resultid="8566" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1276" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7290" />
                    <RANKING order="2" place="2" resultid="7610" />
                    <RANKING order="3" place="3" resultid="8009" />
                    <RANKING order="4" place="4" resultid="7709" />
                    <RANKING order="5" place="5" resultid="8553" />
                    <RANKING order="6" place="6" resultid="8003" />
                    <RANKING order="7" place="7" resultid="7617" />
                    <RANKING order="8" place="8" resultid="8018" />
                    <RANKING order="9" place="9" resultid="8024" />
                    <RANKING order="10" place="10" resultid="9015" />
                    <RANKING order="11" place="-1" resultid="9178" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1277" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7844" />
                    <RANKING order="2" place="2" resultid="7674" />
                    <RANKING order="3" place="3" resultid="8397" />
                    <RANKING order="4" place="4" resultid="7590" />
                    <RANKING order="5" place="5" resultid="8910" />
                    <RANKING order="6" place="6" resultid="8917" />
                    <RANKING order="7" place="7" resultid="7948" />
                    <RANKING order="8" place="8" resultid="7307" />
                    <RANKING order="9" place="-1" resultid="8479" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1278" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7576" />
                    <RANKING order="2" place="2" resultid="8269" />
                    <RANKING order="3" place="3" resultid="7967" />
                    <RANKING order="4" place="-1" resultid="6923" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1279" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6562" />
                    <RANKING order="2" place="2" resultid="7428" />
                    <RANKING order="3" place="3" resultid="6938" />
                    <RANKING order="4" place="4" resultid="6848" />
                    <RANKING order="5" place="5" resultid="7625" />
                    <RANKING order="6" place="6" resultid="7533" />
                    <RANKING order="7" place="-1" resultid="6612" />
                    <RANKING order="8" place="-1" resultid="8675" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1280" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9516" />
                    <RANKING order="2" place="2" resultid="9540" />
                    <RANKING order="3" place="3" resultid="9567" />
                    <RANKING order="4" place="-1" resultid="9602" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10645" daytime="16:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10646" daytime="16:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10647" daytime="16:28" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10648" daytime="16:34" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10649" daytime="16:36" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10650" daytime="16:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10651" daytime="16:44" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10652" daytime="16:48" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1281" daytime="16:52" gender="F" number="38" order="3" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1282" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8153" />
                    <RANKING order="2" place="2" resultid="8147" />
                    <RANKING order="3" place="3" resultid="8358" />
                    <RANKING order="4" place="4" resultid="8264" />
                    <RANKING order="5" place="5" resultid="8207" />
                    <RANKING order="6" place="6" resultid="8318" />
                    <RANKING order="7" place="7" resultid="9270" />
                    <RANKING order="8" place="8" resultid="7135" />
                    <RANKING order="9" place="9" resultid="8739" />
                    <RANKING order="10" place="10" resultid="8258" />
                    <RANKING order="11" place="11" resultid="8594" />
                    <RANKING order="12" place="12" resultid="9607" />
                    <RANKING order="13" place="13" resultid="9022" />
                    <RANKING order="14" place="14" resultid="7161" />
                    <RANKING order="15" place="15" resultid="9414" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1283" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6881" />
                    <RANKING order="2" place="2" resultid="8082" />
                    <RANKING order="3" place="3" resultid="8109" />
                    <RANKING order="4" place="4" resultid="7744" />
                    <RANKING order="5" place="5" resultid="7660" />
                    <RANKING order="6" place="6" resultid="8087" />
                    <RANKING order="7" place="7" resultid="8488" />
                    <RANKING order="8" place="8" resultid="8336" />
                    <RANKING order="9" place="9" resultid="9372" />
                    <RANKING order="10" place="10" resultid="8600" />
                    <RANKING order="11" place="11" resultid="8328" />
                    <RANKING order="12" place="12" resultid="8075" />
                    <RANKING order="13" place="13" resultid="8887" />
                    <RANKING order="14" place="14" resultid="7008" />
                    <RANKING order="15" place="15" resultid="9284" />
                    <RANKING order="16" place="16" resultid="9036" />
                    <RANKING order="17" place="17" resultid="7492" />
                    <RANKING order="18" place="-1" resultid="9157" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1284" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7927" />
                    <RANKING order="2" place="2" resultid="6568" />
                    <RANKING order="3" place="3" resultid="6575" />
                    <RANKING order="4" place="4" resultid="7002" />
                    <RANKING order="5" place="5" resultid="9184" />
                    <RANKING order="6" place="6" resultid="9222" />
                    <RANKING order="7" place="7" resultid="7996" />
                    <RANKING order="8" place="8" resultid="7197" />
                    <RANKING order="9" place="9" resultid="9303" />
                    <RANKING order="10" place="10" resultid="7497" />
                    <RANKING order="11" place="11" resultid="7555" />
                    <RANKING order="12" place="12" resultid="7771" />
                    <RANKING order="13" place="13" resultid="8304" />
                    <RANKING order="14" place="14" resultid="8615" />
                    <RANKING order="15" place="15" resultid="7083" />
                    <RANKING order="16" place="16" resultid="8988" />
                    <RANKING order="17" place="-1" resultid="9589" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1285" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7863" />
                    <RANKING order="2" place="2" resultid="7869" />
                    <RANKING order="3" place="3" resultid="7830" />
                    <RANKING order="4" place="4" resultid="7824" />
                    <RANKING order="5" place="5" resultid="7953" />
                    <RANKING order="6" place="6" resultid="7313" />
                    <RANKING order="7" place="7" resultid="7450" />
                    <RANKING order="8" place="8" resultid="9129" />
                    <RANKING order="9" place="9" resultid="7217" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1286" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8967" />
                    <RANKING order="2" place="2" resultid="7091" />
                    <RANKING order="3" place="3" resultid="9001" />
                    <RANKING order="4" place="4" resultid="7212" />
                    <RANKING order="5" place="5" resultid="7401" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1287" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9087" />
                    <RANKING order="2" place="2" resultid="7568" />
                    <RANKING order="3" place="3" resultid="7336" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1288" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8460" />
                    <RANKING order="2" place="2" resultid="9579" />
                    <RANKING order="3" place="3" resultid="8882" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10653" daytime="16:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10654" daytime="16:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10655" daytime="17:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10656" daytime="17:04" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10657" daytime="17:08" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10658" daytime="17:12" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10659" daytime="17:16" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10660" daytime="17:18" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1289" daytime="17:22" gender="M" number="39" order="4" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1290" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8388" />
                    <RANKING order="2" place="2" resultid="7511" />
                    <RANKING order="3" place="3" resultid="8126" />
                    <RANKING order="4" place="4" resultid="7031" />
                    <RANKING order="5" place="5" resultid="8167" />
                    <RANKING order="6" place="6" resultid="8133" />
                    <RANKING order="7" place="7" resultid="8187" />
                    <RANKING order="8" place="8" resultid="8180" />
                    <RANKING order="9" place="9" resultid="7722" />
                    <RANKING order="10" place="10" resultid="9196" />
                    <RANKING order="11" place="11" resultid="8139" />
                    <RANKING order="12" place="12" resultid="8160" />
                    <RANKING order="13" place="13" resultid="7114" />
                    <RANKING order="14" place="14" resultid="7359" />
                    <RANKING order="15" place="15" resultid="8483" />
                    <RANKING order="16" place="16" resultid="7043" />
                    <RANKING order="17" place="17" resultid="8727" />
                    <RANKING order="18" place="18" resultid="7506" />
                    <RANKING order="19" place="19" resultid="9256" />
                    <RANKING order="20" place="20" resultid="9263" />
                    <RANKING order="21" place="21" resultid="7120" />
                    <RANKING order="22" place="-1" resultid="8233" />
                    <RANKING order="23" place="-1" resultid="8733" />
                    <RANKING order="24" place="-1" resultid="9229" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1291" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7631" />
                    <RANKING order="2" place="2" resultid="8240" />
                    <RANKING order="3" place="3" resultid="8053" />
                    <RANKING order="4" place="4" resultid="7470" />
                    <RANKING order="5" place="5" resultid="8628" />
                    <RANKING order="6" place="6" resultid="6904" />
                    <RANKING order="7" place="7" resultid="8039" />
                    <RANKING order="8" place="8" resultid="8096" />
                    <RANKING order="9" place="9" resultid="8045" />
                    <RANKING order="10" place="10" resultid="8370" />
                    <RANKING order="11" place="11" resultid="9276" />
                    <RANKING order="12" place="12" resultid="9208" />
                    <RANKING order="13" place="13" resultid="9201" />
                    <RANKING order="14" place="14" resultid="7730" />
                    <RANKING order="15" place="15" resultid="7544" />
                    <RANKING order="16" place="16" resultid="8643" />
                    <RANKING order="17" place="17" resultid="7457" />
                    <RANKING order="18" place="18" resultid="8060" />
                    <RANKING order="19" place="19" resultid="6985" />
                    <RANKING order="20" place="20" resultid="8713" />
                    <RANKING order="21" place="21" resultid="7064" />
                    <RANKING order="22" place="22" resultid="6583" />
                    <RANKING order="23" place="23" resultid="7479" />
                    <RANKING order="24" place="24" resultid="7330" />
                    <RANKING order="25" place="25" resultid="7169" />
                    <RANKING order="26" place="26" resultid="7787" />
                    <RANKING order="27" place="27" resultid="9380" />
                    <RANKING order="28" place="28" resultid="8581" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1292" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7905" />
                    <RANKING order="2" place="2" resultid="7611" />
                    <RANKING order="3" place="3" resultid="9326" />
                    <RANKING order="4" place="4" resultid="8004" />
                    <RANKING order="5" place="5" resultid="8311" />
                    <RANKING order="6" place="6" resultid="8010" />
                    <RANKING order="7" place="7" resultid="8032" />
                    <RANKING order="8" place="8" resultid="7464" />
                    <RANKING order="9" place="9" resultid="9149" />
                    <RANKING order="10" place="10" resultid="9250" />
                    <RANKING order="11" place="11" resultid="7977" />
                    <RANKING order="12" place="12" resultid="7778" />
                    <RANKING order="13" place="13" resultid="8949" />
                    <RANKING order="14" place="14" resultid="8019" />
                    <RANKING order="15" place="15" resultid="8025" />
                    <RANKING order="16" place="16" resultid="6968" />
                    <RANKING order="17" place="17" resultid="9420" />
                    <RANKING order="18" place="18" resultid="9460" />
                    <RANKING order="19" place="19" resultid="9446" />
                    <RANKING order="20" place="20" resultid="7342" />
                    <RANKING order="21" place="21" resultid="9425" />
                    <RANKING order="22" place="22" resultid="7794" />
                    <RANKING order="23" place="23" resultid="8807" />
                    <RANKING order="24" place="-1" resultid="7918" />
                    <RANKING order="25" place="-1" resultid="7983" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1293" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6898" />
                    <RANKING order="2" place="2" resultid="6821" />
                    <RANKING order="3" place="3" resultid="7887" />
                    <RANKING order="4" place="4" resultid="7911" />
                    <RANKING order="5" place="5" resultid="8608" />
                    <RANKING order="6" place="6" resultid="7302" />
                    <RANKING order="7" place="7" resultid="6844" />
                    <RANKING order="8" place="8" resultid="9295" />
                    <RANKING order="9" place="9" resultid="8787" />
                    <RANKING order="10" place="10" resultid="9441" />
                    <RANKING order="11" place="11" resultid="9453" />
                    <RANKING order="12" place="12" resultid="8775" />
                    <RANKING order="13" place="13" resultid="8498" />
                    <RANKING order="14" place="-1" resultid="7850" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1294" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8120" />
                    <RANKING order="2" place="2" resultid="6911" />
                    <RANKING order="3" place="3" resultid="9094" />
                    <RANKING order="4" place="4" resultid="8342" />
                    <RANKING order="5" place="5" resultid="7436" />
                    <RANKING order="6" place="6" resultid="9113" />
                    <RANKING order="7" place="7" resultid="7715" />
                    <RANKING order="8" place="8" resultid="9400" />
                    <RANKING order="9" place="9" resultid="7681" />
                    <RANKING order="10" place="10" resultid="8511" />
                    <RANKING order="11" place="11" resultid="6991" />
                    <RANKING order="12" place="12" resultid="9100" />
                    <RANKING order="13" place="13" resultid="8962" />
                    <RANKING order="14" place="14" resultid="7415" />
                    <RANKING order="15" place="15" resultid="7552" />
                    <RANKING order="16" place="16" resultid="9057" />
                    <RANKING order="17" place="17" resultid="7391" />
                    <RANKING order="18" place="-1" resultid="7838" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1295" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7896" />
                    <RANKING order="2" place="2" resultid="8924" />
                    <RANKING order="3" place="3" resultid="7296" />
                    <RANKING order="4" place="4" resultid="9317" />
                    <RANKING order="5" place="5" resultid="8943" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1296" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8352" />
                    <RANKING order="2" place="2" resultid="8408" />
                    <RANKING order="3" place="3" resultid="8365" />
                    <RANKING order="4" place="4" resultid="9121" />
                    <RANKING order="5" place="5" resultid="9547" />
                    <RANKING order="6" place="6" resultid="9572" />
                    <RANKING order="7" place="7" resultid="9386" />
                    <RANKING order="8" place="8" resultid="9559" />
                    <RANKING order="9" place="9" resultid="9584" />
                    <RANKING order="10" place="10" resultid="9510" />
                    <RANKING order="11" place="11" resultid="9595" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10661" daytime="17:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10662" daytime="17:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10663" daytime="17:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10664" daytime="17:36" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10665" daytime="17:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10666" daytime="17:44" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10667" daytime="17:46" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10668" daytime="17:50" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10669" daytime="17:54" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10670" daytime="17:58" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="10671" daytime="18:00" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="10672" daytime="18:04" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="10673" daytime="18:06" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="10674" daytime="18:10" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1297" daytime="18:14" gender="F" number="40" order="5" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1298" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7025" />
                    <RANKING order="2" place="2" resultid="9216" />
                    <RANKING order="3" place="3" resultid="8791" />
                    <RANKING order="4" place="4" resultid="8527" />
                    <RANKING order="5" place="5" resultid="9606" />
                    <RANKING order="6" place="6" resultid="8668" />
                    <RANKING order="7" place="7" resultid="7364" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1299" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6875" />
                    <RANKING order="2" place="2" resultid="7014" />
                    <RANKING order="3" place="3" resultid="7538" />
                    <RANKING order="4" place="3" resultid="8886" />
                    <RANKING order="5" place="5" resultid="9407" />
                    <RANKING order="6" place="6" resultid="9035" />
                    <RANKING order="7" place="7" resultid="7491" />
                    <RANKING order="8" place="8" resultid="9290" />
                    <RANKING order="9" place="9" resultid="8720" />
                    <RANKING order="10" place="10" resultid="7107" />
                    <RANKING order="11" place="11" resultid="9360" />
                    <RANKING order="12" place="-1" resultid="9156" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1300" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7597" />
                    <RANKING order="2" place="2" resultid="7101" />
                    <RANKING order="3" place="3" resultid="7221" />
                    <RANKING order="4" place="4" resultid="7876" />
                    <RANKING order="5" place="5" resultid="6996" />
                    <RANKING order="6" place="6" resultid="8696" />
                    <RANKING order="7" place="7" resultid="8930" />
                    <RANKING order="8" place="8" resultid="9310" />
                    <RANKING order="9" place="9" resultid="6864" />
                    <RANKING order="10" place="10" resultid="9061" />
                    <RANKING order="11" place="11" resultid="8980" />
                    <RANKING order="12" place="12" resultid="8801" />
                    <RANKING order="13" place="13" resultid="7154" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1301" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7283" />
                    <RANKING order="2" place="2" resultid="6830" />
                    <RANKING order="3" place="3" resultid="7320" />
                    <RANKING order="4" place="4" resultid="9067" />
                    <RANKING order="5" place="5" resultid="6840" />
                    <RANKING order="6" place="6" resultid="9128" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1302" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7090" />
                    <RANKING order="2" place="2" resultid="7353" />
                    <RANKING order="3" place="3" resultid="6962" />
                    <RANKING order="4" place="4" resultid="7130" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1303" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7833" />
                    <RANKING order="2" place="2" resultid="6834" />
                    <RANKING order="3" place="3" resultid="9086" />
                    <RANKING order="4" place="4" resultid="9366" />
                    <RANKING order="5" place="5" resultid="7335" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1304" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7406" />
                    <RANKING order="2" place="2" resultid="9529" />
                    <RANKING order="3" place="3" resultid="9505" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10675" daytime="18:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10676" daytime="18:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10677" daytime="18:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10678" daytime="18:22" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10679" daytime="18:24" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10680" daytime="18:26" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1305" daytime="18:28" gender="M" number="41" order="6" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1306" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7036" />
                    <RANKING order="2" place="2" resultid="7149" />
                    <RANKING order="3" place="3" resultid="8586" />
                    <RANKING order="4" place="4" resultid="8955" />
                    <RANKING order="5" place="5" resultid="7174" />
                    <RANKING order="6" place="6" resultid="9344" />
                    <RANKING order="7" place="7" resultid="9262" />
                    <RANKING order="8" place="8" resultid="8663" />
                    <RANKING order="9" place="9" resultid="8795" />
                    <RANKING order="10" place="10" resultid="7054" />
                    <RANKING order="11" place="11" resultid="7113" />
                    <RANKING order="12" place="12" resultid="7255" />
                    <RANKING order="13" place="13" resultid="9437" />
                    <RANKING order="14" place="14" resultid="7505" />
                    <RANKING order="15" place="15" resultid="8764" />
                    <RANKING order="16" place="16" resultid="9333" />
                    <RANKING order="17" place="-1" resultid="8732" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1307" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8627" />
                    <RANKING order="2" place="2" resultid="9141" />
                    <RANKING order="3" place="3" resultid="7143" />
                    <RANKING order="4" place="4" resultid="8688" />
                    <RANKING order="5" place="5" resultid="7232" />
                    <RANKING order="6" place="6" resultid="6856" />
                    <RANKING order="7" place="7" resultid="8102" />
                    <RANKING order="8" place="8" resultid="8642" />
                    <RANKING order="9" place="9" resultid="7478" />
                    <RANKING order="10" place="10" resultid="7241" />
                    <RANKING order="11" place="11" resultid="7168" />
                    <RANKING order="12" place="12" resultid="7249" />
                    <RANKING order="13" place="13" resultid="9353" />
                    <RANKING order="14" place="14" resultid="7227" />
                    <RANKING order="15" place="15" resultid="8709" />
                    <RANKING order="16" place="16" resultid="9379" />
                    <RANKING order="17" place="17" resultid="8770" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1308" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7463" />
                    <RANKING order="2" place="2" resultid="7484" />
                    <RANKING order="3" place="3" resultid="6967" />
                    <RANKING order="4" place="4" resultid="9338" />
                    <RANKING order="5" place="5" resultid="7370" />
                    <RANKING order="6" place="6" resultid="9419" />
                    <RANKING order="7" place="7" resultid="9029" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1309" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7963" />
                    <RANKING order="2" place="1" resultid="8916" />
                    <RANKING order="3" place="3" resultid="8467" />
                    <RANKING order="4" place="4" resultid="6956" />
                    <RANKING order="5" place="5" resultid="8494" />
                    <RANKING order="6" place="6" resultid="7932" />
                    <RANKING order="7" place="7" resultid="8825" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1310" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6950" />
                    <RANKING order="2" place="2" resultid="6910" />
                    <RANKING order="3" place="3" resultid="7414" />
                    <RANKING order="4" place="4" resultid="9093" />
                    <RANKING order="5" place="5" resultid="7347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1311" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8382" />
                    <RANKING order="2" place="2" resultid="8923" />
                    <RANKING order="3" place="3" resultid="8779" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1312" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7202" />
                    <RANKING order="2" place="2" resultid="9116" />
                    <RANKING order="3" place="3" resultid="7192" />
                    <RANKING order="4" place="4" resultid="9321" />
                    <RANKING order="5" place="5" resultid="9120" />
                    <RANKING order="6" place="6" resultid="7409" />
                    <RANKING order="7" place="7" resultid="7421" />
                    <RANKING order="8" place="8" resultid="7796" />
                    <RANKING order="9" place="9" resultid="9523" />
                    <RANKING order="10" place="10" resultid="7208" />
                    <RANKING order="11" place="11" resultid="9553" />
                    <RANKING order="12" place="12" resultid="9509" />
                    <RANKING order="13" place="-1" resultid="9539" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10681" daytime="18:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10682" daytime="18:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10683" daytime="18:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10684" daytime="18:36" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10685" daytime="18:38" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10686" daytime="18:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10687" daytime="18:42" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1313" daytime="18:44" gender="F" number="42" order="7" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1314" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8413" />
                    <RANKING order="2" place="2" resultid="8438" />
                    <RANKING order="3" place="3" resultid="8746" />
                    <RANKING order="4" place="4" resultid="9466" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10688" daytime="18:44" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1315" daytime="18:52" gender="F" number="43" order="8" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1316" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8411" />
                    <RANKING order="2" place="2" resultid="8437" />
                    <RANKING order="3" place="3" resultid="7803" />
                    <RANKING order="4" place="4" resultid="7066" />
                    <RANKING order="5" place="5" resultid="9464" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10689" daytime="18:52" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1317" daytime="18:58" gender="F" number="44" order="9" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1318" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8412" />
                    <RANKING order="2" place="2" resultid="9465" />
                    <RANKING order="3" place="3" resultid="9074" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10690" daytime="18:58" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1319" daytime="19:06" gender="F" number="45" order="10" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1320" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8414" />
                    <RANKING order="2" place="2" resultid="7804" />
                    <RANKING order="3" place="-1" resultid="8439" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10691" daytime="19:06" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1321" daytime="19:12" gender="F" number="46" order="11" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1322" agemax="-1" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7185" />
                    <RANKING order="2" place="2" resultid="9073" />
                    <RANKING order="3" place="3" resultid="9610" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10692" daytime="19:12" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1323" daytime="19:18" gender="M" number="47" order="12" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1324" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8424" />
                    <RANKING order="2" place="2" resultid="7070" />
                    <RANKING order="3" place="3" resultid="8444" />
                    <RANKING order="4" place="4" resultid="7187" />
                    <RANKING order="5" place="5" resultid="8750" />
                    <RANKING order="6" place="6" resultid="9475" />
                    <RANKING order="7" place="7" resultid="8827" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10693" daytime="19:18" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1325" daytime="19:26" gender="M" number="48" order="13" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1326" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7812" />
                    <RANKING order="2" place="2" resultid="9477" />
                    <RANKING order="3" place="3" resultid="8426" />
                    <RANKING order="4" place="4" resultid="8446" />
                    <RANKING order="5" place="5" resultid="7517" />
                    <RANKING order="6" place="6" resultid="8751" />
                    <RANKING order="7" place="7" resultid="7071" />
                    <RANKING order="8" place="8" resultid="7798" />
                    <RANKING order="9" place="9" resultid="9078" />
                    <RANKING order="10" place="10" resultid="9489" />
                    <RANKING order="11" place="11" resultid="7258" />
                    <RANKING order="12" place="-1" resultid="8757" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10694" daytime="19:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10695" daytime="19:32" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1327" daytime="19:40" gender="M" number="49" order="14" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1328" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9488" />
                    <RANKING order="2" place="2" resultid="8425" />
                    <RANKING order="3" place="3" resultid="7811" />
                    <RANKING order="4" place="4" resultid="8445" />
                    <RANKING order="5" place="-1" resultid="9476" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10696" daytime="19:40" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1329" daytime="19:46" gender="M" number="50" order="15" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1330" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8423" />
                    <RANKING order="2" place="2" resultid="8443" />
                    <RANKING order="3" place="3" resultid="7069" />
                    <RANKING order="4" place="4" resultid="9474" />
                    <RANKING order="5" place="5" resultid="8826" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10697" daytime="19:46" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1331" daytime="19:52" gender="M" number="51" order="16" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1332" agemax="-1" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8422" />
                    <RANKING order="2" place="2" resultid="9613" />
                    <RANKING order="3" place="3" resultid="7516" />
                    <RANKING order="4" place="4" resultid="9473" />
                    <RANKING order="5" place="5" resultid="7810" />
                    <RANKING order="6" place="6" resultid="7068" />
                    <RANKING order="7" place="7" resultid="9616" />
                    <RANKING order="8" place="8" resultid="9077" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10698" daytime="19:52" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2025-04-13" daytime="08:55" endtime="13:23" number="5" officialmeeting="08:00" status="OFFICIAL" warmupfrom="07:30" warmupuntil="08:30">
          <EVENTS>
            <EVENT eventid="1333" daytime="08:56" gender="F" number="52" order="1" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1334" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8275" />
                    <RANKING order="2" place="2" resultid="8208" />
                    <RANKING order="3" place="3" resultid="8595" />
                    <RANKING order="4" place="4" resultid="7136" />
                    <RANKING order="5" place="-1" resultid="9271" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1335" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8650" />
                    <RANKING order="2" place="2" resultid="8489" />
                    <RANKING order="3" place="3" resultid="7766" />
                    <RANKING order="4" place="4" resultid="7696" />
                    <RANKING order="5" place="5" resultid="8517" />
                    <RANKING order="6" place="6" resultid="9137" />
                    <RANKING order="7" place="7" resultid="7108" />
                    <RANKING order="8" place="-1" resultid="6809" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1336" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7198" />
                    <RANKING order="2" place="2" resultid="9186" />
                    <RANKING order="3" place="3" resultid="6576" />
                    <RANKING order="4" place="4" resultid="7003" />
                    <RANKING order="5" place="5" resultid="8990" />
                    <RANKING order="6" place="6" resultid="9304" />
                    <RANKING order="7" place="7" resultid="9590" />
                    <RANKING order="8" place="8" resultid="8982" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1337" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7870" />
                    <RANKING order="2" place="2" resultid="7831" />
                    <RANKING order="3" place="3" resultid="7883" />
                    <RANKING order="4" place="4" resultid="8559" />
                    <RANKING order="5" place="5" resultid="6944" />
                    <RANKING order="6" place="6" resultid="7604" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1338" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7647" />
                    <RANKING order="2" place="2" resultid="7402" />
                    <RANKING order="3" place="3" resultid="8904" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1339" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9088" />
                    <RANKING order="2" place="2" resultid="7570" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1340" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="8461" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10699" daytime="08:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10700" daytime="08:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10701" daytime="09:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10702" daytime="09:02" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1341" daytime="09:06" gender="M" number="53" order="2" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1342" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8127" />
                    <RANKING order="2" place="2" resultid="7512" />
                    <RANKING order="3" place="3" resultid="7032" />
                    <RANKING order="4" place="4" resultid="8220" />
                    <RANKING order="5" place="5" resultid="8289" />
                    <RANKING order="6" place="6" resultid="7325" />
                    <RANKING order="7" place="7" resultid="7723" />
                    <RANKING order="8" place="8" resultid="7360" />
                    <RANKING order="9" place="9" resultid="7021" />
                    <RANKING order="10" place="10" resultid="8622" />
                    <RANKING order="11" place="11" resultid="8664" />
                    <RANKING order="12" place="12" resultid="7639" />
                    <RANKING order="13" place="13" resultid="7758" />
                    <RANKING order="14" place="14" resultid="9257" />
                    <RANKING order="15" place="-1" resultid="9346" />
                    <RANKING order="16" place="-1" resultid="6745" />
                    <RANKING order="17" place="-1" resultid="9230" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1343" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9277" />
                    <RANKING order="2" place="2" resultid="7471" />
                    <RANKING order="3" place="3" resultid="7632" />
                    <RANKING order="4" place="4" resultid="9143" />
                    <RANKING order="5" place="5" resultid="8629" />
                    <RANKING order="6" place="6" resultid="8637" />
                    <RANKING order="7" place="7" resultid="6905" />
                    <RANKING order="8" place="8" resultid="9202" />
                    <RANKING order="9" place="9" resultid="7667" />
                    <RANKING order="10" place="10" resultid="8046" />
                    <RANKING order="11" place="11" resultid="7752" />
                    <RANKING order="12" place="12" resultid="8567" />
                    <RANKING order="13" place="13" resultid="8297" />
                    <RANKING order="14" place="14" resultid="7688" />
                    <RANKING order="15" place="15" resultid="8704" />
                    <RANKING order="16" place="16" resultid="7237" />
                    <RANKING order="17" place="17" resultid="6889" />
                    <RANKING order="18" place="18" resultid="8995" />
                    <RANKING order="19" place="19" resultid="6974" />
                    <RANKING order="20" place="-1" resultid="8116" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1344" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7291" />
                    <RANKING order="2" place="2" resultid="9150" />
                    <RANKING order="3" place="3" resultid="7485" />
                    <RANKING order="4" place="4" resultid="7779" />
                    <RANKING order="5" place="5" resultid="9016" />
                    <RANKING order="6" place="6" resultid="8532" />
                    <RANKING order="7" place="7" resultid="7618" />
                    <RANKING order="8" place="8" resultid="9339" />
                    <RANKING order="9" place="9" resultid="9030" />
                    <RANKING order="10" place="-1" resultid="6682" />
                    <RANKING order="11" place="-1" resultid="9179" />
                    <RANKING order="12" place="-1" resultid="8026" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1345" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6899" />
                    <RANKING order="2" place="2" resultid="7675" />
                    <RANKING order="3" place="3" resultid="8348" />
                    <RANKING order="4" place="4" resultid="8377" />
                    <RANKING order="5" place="5" resultid="6957" />
                    <RANKING order="6" place="6" resultid="7308" />
                    <RANKING order="7" place="7" resultid="6918" />
                    <RANKING order="8" place="8" resultid="9296" />
                    <RANKING order="9" place="-1" resultid="7958" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1346" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7577" />
                    <RANKING order="2" place="2" resultid="7716" />
                    <RANKING order="3" place="3" resultid="9095" />
                    <RANKING order="4" place="4" resultid="9401" />
                    <RANKING order="5" place="5" resultid="6992" />
                    <RANKING order="6" place="-1" resultid="7387" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1347" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7429" />
                    <RANKING order="2" place="2" resultid="8894" />
                    <RANKING order="3" place="3" resultid="6939" />
                    <RANKING order="4" place="4" resultid="6849" />
                    <RANKING order="5" place="5" resultid="7297" />
                    <RANKING order="6" place="6" resultid="7443" />
                    <RANKING order="7" place="7" resultid="8676" />
                    <RANKING order="8" place="8" resultid="7534" />
                    <RANKING order="9" place="-1" resultid="6563" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1348" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7203" />
                    <RANKING order="2" place="2" resultid="9189" />
                    <RANKING order="3" place="3" resultid="9573" />
                    <RANKING order="4" place="4" resultid="9122" />
                    <RANKING order="5" place="5" resultid="7422" />
                    <RANKING order="6" place="6" resultid="9548" />
                    <RANKING order="7" place="7" resultid="9541" />
                    <RANKING order="8" place="8" resultid="9554" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10703" daytime="09:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10704" daytime="09:08" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10705" daytime="09:12" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10706" daytime="09:14" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10707" daytime="09:16" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10708" daytime="09:18" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10709" daytime="09:20" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10710" daytime="09:22" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10711" daytime="09:26" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1349" daytime="09:28" gender="F" number="54" order="3" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1350" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8154" />
                    <RANKING order="2" place="2" resultid="8201" />
                    <RANKING order="3" place="3" resultid="8148" />
                    <RANKING order="4" place="4" resultid="8265" />
                    <RANKING order="5" place="5" resultid="8359" />
                    <RANKING order="6" place="6" resultid="8319" />
                    <RANKING order="7" place="7" resultid="9050" />
                    <RANKING order="8" place="8" resultid="8740" />
                    <RANKING order="9" place="9" resultid="9023" />
                    <RANKING order="10" place="10" resultid="8657" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1351" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8110" />
                    <RANKING order="2" place="2" resultid="7661" />
                    <RANKING order="3" place="3" resultid="8088" />
                    <RANKING order="4" place="4" resultid="8601" />
                    <RANKING order="5" place="5" resultid="8649" />
                    <RANKING order="6" place="6" resultid="7745" />
                    <RANKING order="7" place="7" resultid="9373" />
                    <RANKING order="8" place="8" resultid="8888" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1352" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6569" />
                    <RANKING order="2" place="2" resultid="7928" />
                    <RANKING order="3" place="3" resultid="7703" />
                    <RANKING order="4" place="4" resultid="7997" />
                    <RANKING order="5" place="5" resultid="8932" />
                    <RANKING order="6" place="6" resultid="9185" />
                    <RANKING order="7" place="7" resultid="7498" />
                    <RANKING order="8" place="8" resultid="9223" />
                    <RANKING order="9" place="9" resultid="9237" />
                    <RANKING order="10" place="10" resultid="7772" />
                    <RANKING order="11" place="11" resultid="7084" />
                    <RANKING order="12" place="12" resultid="8616" />
                    <RANKING order="13" place="13" resultid="8989" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1353" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7864" />
                    <RANKING order="2" place="2" resultid="7825" />
                    <RANKING order="3" place="3" resultid="7451" />
                    <RANKING order="4" place="4" resultid="7528" />
                    <RANKING order="5" place="-1" resultid="6648" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1354" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8968" />
                    <RANKING order="2" place="2" resultid="7213" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1355" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7569" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1356" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9535" />
                    <RANKING order="2" place="2" resultid="9580" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10712" daytime="09:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10713" daytime="09:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10714" daytime="09:42" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10715" daytime="09:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10716" daytime="09:54" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1357" daytime="10:02" gender="M" number="55" order="4" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1358" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7038" />
                    <RANKING order="2" place="2" resultid="7724" />
                    <RANKING order="3" place="3" resultid="8140" />
                    <RANKING order="4" place="4" resultid="8623" />
                    <RANKING order="5" place="5" resultid="7044" />
                    <RANKING order="6" place="6" resultid="8175" />
                    <RANKING order="7" place="-1" resultid="7513" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1359" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8054" />
                    <RANKING order="2" place="2" resultid="8241" />
                    <RANKING order="3" place="3" resultid="8040" />
                    <RANKING order="4" place="4" resultid="7654" />
                    <RANKING order="5" place="5" resultid="9203" />
                    <RANKING order="6" place="6" resultid="8047" />
                    <RANKING order="7" place="7" resultid="8975" />
                    <RANKING order="8" place="8" resultid="8371" />
                    <RANKING order="9" place="9" resultid="9209" />
                    <RANKING order="10" place="10" resultid="7668" />
                    <RANKING order="11" place="11" resultid="8283" />
                    <RANKING order="12" place="12" resultid="9278" />
                    <RANKING order="13" place="13" resultid="8473" />
                    <RANKING order="14" place="14" resultid="8061" />
                    <RANKING order="15" place="15" resultid="6986" />
                    <RANKING order="16" place="16" resultid="6584" />
                    <RANKING order="17" place="17" resultid="7065" />
                    <RANKING order="18" place="-1" resultid="7545" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1360" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7906" />
                    <RANKING order="2" place="2" resultid="8033" />
                    <RANKING order="3" place="3" resultid="9327" />
                    <RANKING order="4" place="4" resultid="8011" />
                    <RANKING order="5" place="5" resultid="7710" />
                    <RANKING order="6" place="6" resultid="8939" />
                    <RANKING order="7" place="7" resultid="8312" />
                    <RANKING order="8" place="8" resultid="9151" />
                    <RANKING order="9" place="9" resultid="7780" />
                    <RANKING order="10" place="10" resultid="9251" />
                    <RANKING order="11" place="11" resultid="7619" />
                    <RANKING order="12" place="12" resultid="9447" />
                    <RANKING order="13" place="13" resultid="9461" />
                    <RANKING order="14" place="-1" resultid="7919" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1361" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6822" />
                    <RANKING order="2" place="2" resultid="7888" />
                    <RANKING order="3" place="3" resultid="8911" />
                    <RANKING order="4" place="4" resultid="7591" />
                    <RANKING order="5" place="5" resultid="6845" />
                    <RANKING order="6" place="6" resultid="9297" />
                    <RANKING order="7" place="7" resultid="6980" />
                    <RANKING order="8" place="8" resultid="9454" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1362" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8121" />
                    <RANKING order="2" place="2" resultid="7437" />
                    <RANKING order="3" place="3" resultid="7717" />
                    <RANKING order="4" place="4" resultid="9114" />
                    <RANKING order="5" place="5" resultid="6924" />
                    <RANKING order="6" place="6" resultid="7682" />
                    <RANKING order="7" place="7" resultid="9101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1363" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7858" />
                    <RANKING order="2" place="2" resultid="7897" />
                    <RANKING order="3" place="3" resultid="8925" />
                    <RANKING order="4" place="4" resultid="8944" />
                    <RANKING order="5" place="5" resultid="7444" />
                    <RANKING order="6" place="6" resultid="9318" />
                    <RANKING order="7" place="7" resultid="7626" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1364" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9387" />
                    <RANKING order="2" place="2" resultid="9568" />
                    <RANKING order="3" place="3" resultid="9560" />
                    <RANKING order="4" place="4" resultid="9596" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10717" daytime="10:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10718" daytime="10:08" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10719" daytime="10:16" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10720" daytime="10:24" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10721" daytime="10:30" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10722" daytime="10:36" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10723" daytime="10:42" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10724" daytime="10:48" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1365" daytime="10:54" gender="F" number="56" order="5" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1366" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8276" />
                    <RANKING order="2" place="2" resultid="8155" />
                    <RANKING order="3" place="3" resultid="8320" />
                    <RANKING order="4" place="4" resultid="8259" />
                    <RANKING order="5" place="5" resultid="9432" />
                    <RANKING order="6" place="6" resultid="7026" />
                    <RANKING order="7" place="7" resultid="7137" />
                    <RANKING order="8" place="8" resultid="9608" />
                    <RANKING order="9" place="9" resultid="7738" />
                    <RANKING order="10" place="10" resultid="8195" />
                    <RANKING order="11" place="11" resultid="8792" />
                    <RANKING order="12" place="12" resultid="8528" />
                    <RANKING order="13" place="13" resultid="7162" />
                    <RANKING order="14" place="14" resultid="8669" />
                    <RANKING order="15" place="15" resultid="7365" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1367" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8248" />
                    <RANKING order="2" place="2" resultid="8329" />
                    <RANKING order="3" place="3" resultid="6882" />
                    <RANKING order="4" place="4" resultid="8089" />
                    <RANKING order="5" place="5" resultid="6876" />
                    <RANKING order="6" place="6" resultid="8602" />
                    <RANKING order="7" place="7" resultid="7015" />
                    <RANKING order="8" place="8" resultid="8889" />
                    <RANKING order="9" place="9" resultid="7540" />
                    <RANKING order="10" place="10" resultid="7009" />
                    <RANKING order="11" place="11" resultid="9285" />
                    <RANKING order="12" place="12" resultid="9037" />
                    <RANKING order="13" place="13" resultid="9408" />
                    <RANKING order="14" place="14" resultid="8721" />
                    <RANKING order="15" place="-1" resultid="9158" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1368" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7598" />
                    <RANKING order="2" place="2" resultid="6577" />
                    <RANKING order="3" place="3" resultid="6570" />
                    <RANKING order="4" place="4" resultid="7102" />
                    <RANKING order="5" place="5" resultid="7991" />
                    <RANKING order="6" place="6" resultid="7222" />
                    <RANKING order="7" place="7" resultid="7998" />
                    <RANKING order="8" place="8" resultid="6997" />
                    <RANKING order="9" place="9" resultid="8697" />
                    <RANKING order="10" place="10" resultid="7773" />
                    <RANKING order="11" place="11" resultid="9311" />
                    <RANKING order="12" place="12" resultid="7085" />
                    <RANKING order="13" place="13" resultid="9062" />
                    <RANKING order="14" place="14" resultid="8983" />
                    <RANKING order="15" place="15" resultid="7155" />
                    <RANKING order="16" place="-1" resultid="7499" />
                    <RANKING order="17" place="-1" resultid="8802" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1369" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7285" />
                    <RANKING order="2" place="2" resultid="6831" />
                    <RANKING order="3" place="3" resultid="8560" />
                    <RANKING order="4" place="4" resultid="7605" />
                    <RANKING order="5" place="5" resultid="7938" />
                    <RANKING order="6" place="6" resultid="7314" />
                    <RANKING order="7" place="7" resultid="9130" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1370" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7092" />
                    <RANKING order="2" place="2" resultid="8969" />
                    <RANKING order="3" place="3" resultid="7403" />
                    <RANKING order="4" place="4" resultid="9002" />
                    <RANKING order="5" place="5" resultid="7354" />
                    <RANKING order="6" place="6" resultid="6963" />
                    <RANKING order="7" place="7" resultid="7131" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1371" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7834" />
                    <RANKING order="2" place="2" resultid="6835" />
                    <RANKING order="3" place="3" resultid="8683" />
                    <RANKING order="4" place="4" resultid="7337" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1372" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7584" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10725" daytime="10:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10726" daytime="10:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10727" daytime="11:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10728" daytime="11:04" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10729" daytime="11:08" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10730" daytime="11:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10731" daytime="11:14" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10732" daytime="11:16" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1373" daytime="11:18" gender="M" number="57" order="6" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1374" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8389" />
                    <RANKING order="2" place="2" resultid="8128" />
                    <RANKING order="3" place="3" resultid="8588" />
                    <RANKING order="4" place="4" resultid="8188" />
                    <RANKING order="5" place="5" resultid="7175" />
                    <RANKING order="6" place="6" resultid="7150" />
                    <RANKING order="7" place="7" resultid="8134" />
                    <RANKING order="8" place="8" resultid="8957" />
                    <RANKING order="9" place="9" resultid="8181" />
                    <RANKING order="10" place="10" resultid="8168" />
                    <RANKING order="11" place="11" resultid="8797" />
                    <RANKING order="12" place="12" resultid="8161" />
                    <RANKING order="13" place="13" resultid="8234" />
                    <RANKING order="14" place="14" resultid="9264" />
                    <RANKING order="15" place="15" resultid="7640" />
                    <RANKING order="16" place="16" resultid="8214" />
                    <RANKING order="17" place="17" resultid="7256" />
                    <RANKING order="18" place="18" resultid="8141" />
                    <RANKING order="19" place="19" resultid="7055" />
                    <RANKING order="20" place="20" resultid="7759" />
                    <RANKING order="21" place="21" resultid="8765" />
                    <RANKING order="22" place="22" resultid="8821" />
                    <RANKING order="23" place="-1" resultid="8734" />
                    <RANKING order="24" place="-1" resultid="6746" />
                    <RANKING order="25" place="-1" resultid="9347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1375" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7633" />
                    <RANKING order="2" place="2" resultid="8630" />
                    <RANKING order="3" place="3" resultid="9144" />
                    <RANKING order="4" place="4" resultid="7144" />
                    <RANKING order="5" place="5" resultid="8690" />
                    <RANKING order="6" place="6" resultid="8117" />
                    <RANKING order="7" place="7" resultid="7472" />
                    <RANKING order="8" place="8" resultid="8103" />
                    <RANKING order="9" place="9" resultid="8644" />
                    <RANKING order="10" place="10" resultid="8976" />
                    <RANKING order="11" place="11" resultid="7731" />
                    <RANKING order="12" place="12" resultid="8714" />
                    <RANKING order="13" place="13" resultid="8372" />
                    <RANKING order="14" place="14" resultid="7458" />
                    <RANKING order="15" place="15" resultid="7689" />
                    <RANKING order="16" place="16" resultid="7242" />
                    <RANKING order="17" place="17" resultid="9354" />
                    <RANKING order="18" place="18" resultid="8811" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1376" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7292" />
                    <RANKING order="2" place="2" resultid="7612" />
                    <RANKING order="3" place="3" resultid="7465" />
                    <RANKING order="4" place="4" resultid="7486" />
                    <RANKING order="5" place="5" resultid="8005" />
                    <RANKING order="6" place="6" resultid="8012" />
                    <RANKING order="7" place="7" resultid="8313" />
                    <RANKING order="8" place="8" resultid="8950" />
                    <RANKING order="9" place="9" resultid="9340" />
                    <RANKING order="10" place="10" resultid="6969" />
                    <RANKING order="11" place="11" resultid="7907" />
                    <RANKING order="12" place="12" resultid="7371" />
                    <RANKING order="13" place="-1" resultid="7984" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1377" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7912" />
                    <RANKING order="2" place="2" resultid="7845" />
                    <RANKING order="3" place="3" resultid="7964" />
                    <RANKING order="4" place="4" resultid="8398" />
                    <RANKING order="5" place="5" resultid="8918" />
                    <RANKING order="6" place="6" resultid="8609" />
                    <RANKING order="7" place="7" resultid="8468" />
                    <RANKING order="8" place="-1" resultid="7933" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1378" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7968" />
                    <RANKING order="2" place="2" resultid="8343" />
                    <RANKING order="3" place="3" resultid="6951" />
                    <RANKING order="4" place="4" resultid="6912" />
                    <RANKING order="5" place="5" resultid="7416" />
                    <RANKING order="6" place="6" resultid="7348" />
                    <RANKING order="7" place="-1" resultid="7839" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1379" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8383" />
                    <RANKING order="2" place="2" resultid="7430" />
                    <RANKING order="3" place="3" resultid="8780" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1380" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9517" />
                    <RANKING order="2" place="2" resultid="9123" />
                    <RANKING order="3" place="3" resultid="9117" />
                    <RANKING order="4" place="4" resultid="7423" />
                    <RANKING order="5" place="5" resultid="7797" />
                    <RANKING order="6" place="6" resultid="9542" />
                    <RANKING order="7" place="7" resultid="7193" />
                    <RANKING order="8" place="8" resultid="9499" />
                    <RANKING order="9" place="9" resultid="9561" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10733" daytime="11:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10734" daytime="11:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10735" daytime="11:26" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10736" daytime="11:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10737" daytime="11:32" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10738" daytime="11:36" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10739" daytime="11:38" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10740" daytime="11:42" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10741" daytime="11:44" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10742" daytime="11:48" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1381" daytime="11:50" gender="F" number="58" order="7" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1382" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8415" />
                    <RANKING order="2" place="2" resultid="8440" />
                    <RANKING order="3" place="3" resultid="9467" />
                    <RANKING order="4" place="4" resultid="8747" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10743" daytime="11:50" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1383" daytime="11:58" gender="F" number="59" order="8" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1384" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8418" />
                    <RANKING order="2" place="2" resultid="8442" />
                    <RANKING order="3" place="3" resultid="7806" />
                    <RANKING order="4" place="4" resultid="7067" />
                    <RANKING order="5" place="5" resultid="9469" />
                    <RANKING order="6" place="6" resultid="8748" />
                    <RANKING order="7" place="7" resultid="9076" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10744" daytime="11:58" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1385" daytime="12:04" gender="F" number="60" order="9" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1386" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8417" />
                    <RANKING order="2" place="2" resultid="9468" />
                    <RANKING order="3" place="3" resultid="9075" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10745" daytime="12:04" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1387" daytime="12:10" gender="F" number="61" order="10" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1388" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8416" />
                    <RANKING order="2" place="2" resultid="8441" />
                    <RANKING order="3" place="3" resultid="7805" />
                    <RANKING order="4" place="4" resultid="6890" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10746" daytime="12:10" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1389" daytime="12:16" gender="F" number="62" order="11" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1390" agemax="-1" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="7186" />
                    <RANKING order="2" place="2" resultid="9611" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10747" daytime="12:16" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1391" daytime="12:22" gender="M" number="63" order="12" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1392" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8431" />
                    <RANKING order="2" place="2" resultid="7075" />
                    <RANKING order="3" place="3" resultid="8450" />
                    <RANKING order="4" place="4" resultid="7188" />
                    <RANKING order="5" place="5" resultid="8753" />
                    <RANKING order="6" place="6" resultid="8829" />
                    <RANKING order="7" place="-1" resultid="9482" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10748" daytime="12:22" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1393" daytime="12:28" gender="M" number="64" order="13" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1394" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8430" />
                    <RANKING order="2" place="2" resultid="7815" />
                    <RANKING order="3" place="3" resultid="9481" />
                    <RANKING order="4" place="4" resultid="8449" />
                    <RANKING order="5" place="5" resultid="7074" />
                    <RANKING order="6" place="6" resultid="8752" />
                    <RANKING order="7" place="7" resultid="7519" />
                    <RANKING order="8" place="8" resultid="9491" />
                    <RANKING order="9" place="9" resultid="7799" />
                    <RANKING order="10" place="10" resultid="7259" />
                    <RANKING order="11" place="11" resultid="7394" />
                    <RANKING order="12" place="12" resultid="8758" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10749" daytime="12:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10750" daytime="12:34" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1395" daytime="12:40" gender="M" number="65" order="14" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1396" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8429" />
                    <RANKING order="2" place="2" resultid="9480" />
                    <RANKING order="3" place="3" resultid="7814" />
                    <RANKING order="4" place="4" resultid="8448" />
                    <RANKING order="5" place="5" resultid="9080" />
                    <RANKING order="6" place="6" resultid="9490" />
                    <RANKING order="7" place="-1" resultid="7393" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10751" daytime="12:40" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1397" daytime="12:46" gender="M" number="66" order="15" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1398" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8428" />
                    <RANKING order="2" place="2" resultid="8447" />
                    <RANKING order="3" place="3" resultid="7073" />
                    <RANKING order="4" place="-1" resultid="8828" />
                    <RANKING order="5" place="-1" resultid="9479" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10752" daytime="12:46" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1399" daytime="12:52" gender="M" number="67" order="16" round="TIM" status="OFFICIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1400" agemax="-1" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="8427" />
                    <RANKING order="2" place="2" resultid="9478" />
                    <RANKING order="3" place="3" resultid="9614" />
                    <RANKING order="4" place="4" resultid="7518" />
                    <RANKING order="5" place="5" resultid="7072" />
                    <RANKING order="6" place="6" resultid="7813" />
                    <RANKING order="7" place="7" resultid="9617" />
                    <RANKING order="8" place="8" resultid="9079" />
                    <RANKING order="9" place="9" resultid="7392" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10753" daytime="12:52" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="13038" nation="BRA" region="PR" clubid="7079" swrid="93759" name="Associação De Pais E Atletas De Natação Ws/Crb" shortname="Apan/Ws">
          <ATHLETES>
            <ATHLETE firstname="Manuela" lastname="Cravcenco Marcondes" birthdate="2012-06-23" gender="F" nation="BRA" license="406866" swrid="5725987" athleteid="7156" externalid="406866">
              <RESULTS>
                <RESULT eventid="1095" points="147" swimtime="00:00:46.21" resultid="7157" heatid="10495" lane="3" entrytime="00:00:45.42" entrycourse="LCM" />
                <RESULT eventid="1179" points="223" swimtime="00:00:48.05" resultid="7158" heatid="10562" lane="8" entrytime="00:00:47.73" entrycourse="LCM" />
                <RESULT eventid="1147" points="274" swimtime="00:01:19.56" resultid="7159" heatid="10526" lane="8" entrytime="00:01:20.83" entrycourse="LCM" />
                <RESULT eventid="1227" points="300" swimtime="00:00:35.23" resultid="7160" heatid="10602" lane="3" entrytime="00:00:35.38" entrycourse="LCM" />
                <RESULT eventid="1281" points="251" swimtime="00:02:57.87" resultid="7161" heatid="10654" lane="1" entrytime="00:03:15.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                    <SPLIT distance="100" swimtime="00:01:22.66" />
                    <SPLIT distance="150" swimtime="00:02:11.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="240" swimtime="00:01:31.86" resultid="7162" heatid="10727" lane="0" entrytime="00:01:38.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Ferreira" birthdate="2012-12-29" gender="F" nation="BRA" license="382235" swrid="5602538" athleteid="7132" externalid="382235">
              <RESULTS>
                <RESULT eventid="1147" points="387" swimtime="00:01:10.91" resultid="7133" heatid="10526" lane="3" entrytime="00:01:19.54" entrycourse="LCM" />
                <RESULT eventid="1227" points="388" swimtime="00:00:32.35" resultid="7134" heatid="10604" lane="0" entrytime="00:00:32.45" entrycourse="LCM" />
                <RESULT eventid="1281" points="383" swimtime="00:02:34.46" resultid="7135" heatid="10655" lane="4" entrytime="00:02:36.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                    <SPLIT distance="100" swimtime="00:01:13.57" />
                    <SPLIT distance="150" swimtime="00:01:55.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="286" swimtime="00:01:23.75" resultid="7136" heatid="10700" lane="3" entrytime="00:01:26.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="293" swimtime="00:01:25.95" resultid="7137" heatid="10728" lane="1" entrytime="00:01:28.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Daniele Silva" birthdate="2010-07-06" gender="F" nation="BRA" license="359593" swrid="5588628" athleteid="7097" externalid="359593" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1063" points="362" swimtime="00:02:52.63" resultid="7098" heatid="10471" lane="8" entrytime="00:02:54.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.68" />
                    <SPLIT distance="100" swimtime="00:01:21.75" />
                    <SPLIT distance="150" swimtime="00:02:07.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="445" swimtime="00:01:07.69" resultid="7099" heatid="10532" lane="2" entrytime="00:01:05.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="487" swimtime="00:00:30.00" resultid="7100" heatid="10609" lane="8" entrytime="00:00:29.13" entrycourse="LCM" />
                <RESULT eventid="1297" points="446" swimtime="00:00:35.14" resultid="7101" heatid="10680" lane="2" entrytime="00:00:34.55" entrycourse="LCM" />
                <RESULT eventid="1365" points="392" swimtime="00:01:18.03" resultid="7102" heatid="10731" lane="2" entrytime="00:01:16.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Cravcenco Marcondes" birthdate="2011-05-06" gender="M" nation="BRA" license="406867" swrid="5723023" athleteid="7163" externalid="406867">
              <RESULTS>
                <RESULT eventid="1103" points="288" swimtime="00:00:33.71" resultid="7164" heatid="10503" lane="6" entrytime="00:00:35.47" entrycourse="LCM" />
                <RESULT eventid="1187" points="188" swimtime="00:00:45.28" resultid="7165" heatid="10570" lane="5" entrytime="00:00:45.81" entrycourse="LCM" />
                <RESULT eventid="1155" points="288" swimtime="00:01:10.22" resultid="7166" heatid="10541" lane="6" entrytime="00:01:10.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="325" swimtime="00:00:30.41" resultid="7167" heatid="10618" lane="5" entrytime="00:00:30.30" entrycourse="LCM" />
                <RESULT eventid="1305" points="229" swimtime="00:00:38.47" resultid="7168" heatid="10684" lane="6" entrytime="00:00:38.42" entrycourse="LCM" />
                <RESULT eventid="1289" points="254" swimtime="00:02:40.98" resultid="7169" heatid="10665" lane="5" entrytime="00:02:42.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                    <SPLIT distance="100" swimtime="00:01:15.48" />
                    <SPLIT distance="150" swimtime="00:01:59.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Da Reginalda" birthdate="2012-11-09" gender="M" nation="BRA" license="400275" swrid="5717253" athleteid="7145" externalid="400275">
              <RESULTS>
                <RESULT eventid="1071" points="313" swimtime="00:02:44.69" resultid="7146" heatid="10475" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                    <SPLIT distance="100" swimtime="00:01:21.39" />
                    <SPLIT distance="150" swimtime="00:02:06.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="358" swimtime="00:01:05.31" resultid="7147" heatid="10543" lane="5" entrytime="00:01:06.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="383" swimtime="00:00:28.79" resultid="7148" heatid="10620" lane="1" entrytime="00:00:29.43" entrycourse="LCM" />
                <RESULT eventid="1305" points="329" swimtime="00:00:34.11" resultid="7149" heatid="10685" lane="8" entrytime="00:00:35.44" entrycourse="LCM" />
                <RESULT eventid="1373" points="308" swimtime="00:01:16.39" resultid="7150" heatid="10738" lane="0" entrytime="00:01:15.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Reis" birthdate="2008-04-07" gender="F" nation="BRA" license="378820" swrid="5600243" athleteid="7126" externalid="378820" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1095" points="201" swimtime="00:00:41.65" resultid="7127" heatid="10496" lane="9" entrytime="00:00:42.43" entrycourse="LCM" />
                <RESULT eventid="1147" points="281" swimtime="00:01:18.92" resultid="7128" heatid="10526" lane="6" entrytime="00:01:19.75" entrycourse="LCM" />
                <RESULT eventid="1227" points="266" swimtime="00:00:36.70" resultid="7129" heatid="10603" lane="9" entrytime="00:00:34.93" entrycourse="LCM" />
                <RESULT eventid="1297" points="248" swimtime="00:00:42.74" resultid="7130" heatid="10678" lane="7" entrytime="00:00:42.05" entrycourse="LCM" />
                <RESULT eventid="1365" points="228" swimtime="00:01:33.46" resultid="7131" heatid="10727" lane="4" entrytime="00:01:30.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Ueda Pritzsche" birthdate="2012-02-07" gender="M" nation="BRA" license="417110" swrid="5756912" athleteid="7170" externalid="417110">
              <RESULTS>
                <RESULT eventid="1103" points="255" swimtime="00:00:35.09" resultid="7171" heatid="10504" lane="0" entrytime="00:00:34.61" entrycourse="LCM" />
                <RESULT eventid="1155" points="277" swimtime="00:01:11.10" resultid="7172" heatid="10540" lane="1" entrytime="00:01:13.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="321" swimtime="00:00:30.51" resultid="7173" heatid="10617" lane="4" entrytime="00:00:30.98" entrycourse="LCM" />
                <RESULT eventid="1305" points="284" swimtime="00:00:35.81" resultid="7174" heatid="10684" lane="1" entrytime="00:00:40.28" entrycourse="LCM" />
                <RESULT eventid="1373" points="312" swimtime="00:01:16.05" resultid="7175" heatid="10737" lane="1" entrytime="00:01:18.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Rosa Silva" birthdate="2011-03-25" gender="F" nation="BRA" license="392120" swrid="5602579" athleteid="7121" externalid="392120">
              <RESULTS>
                <RESULT eventid="1095" points="186" swimtime="00:00:42.73" resultid="7122" heatid="10494" lane="0" />
                <RESULT eventid="1179" points="223" swimtime="00:00:48.02" resultid="7123" heatid="10562" lane="2" entrytime="00:00:45.19" entrycourse="LCM" />
                <RESULT eventid="1147" points="292" swimtime="00:01:17.92" resultid="7124" heatid="10526" lane="4" entrytime="00:01:18.79" entrycourse="LCM" />
                <RESULT eventid="1265" points="250" swimtime="00:03:20.00" resultid="7125" heatid="10640" lane="0" entrytime="00:03:27.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.95" />
                    <SPLIT distance="100" swimtime="00:01:37.59" />
                    <SPLIT distance="150" swimtime="00:02:35.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Bernardi Iurk" birthdate="2012-04-14" gender="M" nation="BRA" license="406940" swrid="5717245" athleteid="7109" externalid="406940">
              <RESULTS>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 11:15)" eventid="1103" status="DSQ" swimtime="00:00:36.15" resultid="7110" heatid="10502" lane="5" entrytime="00:00:39.97" entrycourse="LCM" />
                <RESULT eventid="1155" points="290" swimtime="00:01:10.08" resultid="7111" heatid="10542" lane="7" entrytime="00:01:09.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="309" swimtime="00:00:30.91" resultid="7112" heatid="10617" lane="6" entrytime="00:00:31.09" entrycourse="LCM" />
                <RESULT eventid="1305" points="173" swimtime="00:00:42.19" resultid="7113" heatid="10684" lane="0" entrytime="00:00:41.80" entrycourse="LCM" />
                <RESULT eventid="1289" points="269" swimtime="00:02:37.87" resultid="7114" heatid="10665" lane="6" entrytime="00:02:44.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                    <SPLIT distance="100" swimtime="00:01:15.97" />
                    <SPLIT distance="150" swimtime="00:01:58.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Da Costa Riekes" birthdate="2008-06-19" gender="F" nation="BRA" license="331686" swrid="5600143" athleteid="7086" externalid="331686" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1095" points="414" swimtime="00:00:32.76" resultid="7087" heatid="10498" lane="2" entrytime="00:00:31.38" entrycourse="LCM" />
                <RESULT eventid="1147" points="565" swimtime="00:01:02.52" resultid="7088" heatid="10534" lane="2" entrytime="00:01:02.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="544" swimtime="00:00:28.91" resultid="7089" heatid="10609" lane="2" entrytime="00:00:28.82" entrycourse="LCM" />
                <RESULT eventid="1297" points="461" swimtime="00:00:34.75" resultid="7090" heatid="10680" lane="8" entrytime="00:00:35.66" entrycourse="LCM" />
                <RESULT eventid="1281" points="502" swimtime="00:02:21.12" resultid="7091" heatid="10660" lane="8" entrytime="00:02:19.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.15" />
                    <SPLIT distance="100" swimtime="00:01:06.79" />
                    <SPLIT distance="150" swimtime="00:01:44.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="431" swimtime="00:01:15.62" resultid="7092" heatid="10732" lane="0" entrytime="00:01:13.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Lima Andrade" birthdate="2007-02-09" gender="F" nation="BRA" license="329417" swrid="5820330" athleteid="7176" externalid="329417">
              <RESULTS>
                <RESULT eventid="1095" points="494" swimtime="00:00:30.89" resultid="7177" heatid="10498" lane="5" entrytime="00:00:30.22" entrycourse="LCM" />
                <RESULT eventid="1079" points="418" swimtime="00:03:03.82" resultid="7178" heatid="10485" lane="5" entrytime="00:02:56.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                    <SPLIT distance="100" swimtime="00:01:25.81" />
                    <SPLIT distance="150" swimtime="00:02:14.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="504" swimtime="00:00:36.62" resultid="7179" heatid="10565" lane="4" entrytime="00:00:35.02" entrycourse="LCM" />
                <RESULT eventid="1211" points="463" swimtime="00:01:22.88" resultid="7180" heatid="10589" lane="2" entrytime="00:01:18.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="478" swimtime="00:02:41.20" resultid="7181" heatid="10644" lane="6" entrytime="00:02:38.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                    <SPLIT distance="100" swimtime="00:01:17.15" />
                    <SPLIT distance="150" swimtime="00:02:02.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Sieck" birthdate="2011-01-20" gender="F" nation="BRA" license="382234" swrid="5602584" athleteid="7103" externalid="382234">
              <RESULTS>
                <RESULT eventid="1095" points="215" swimtime="00:00:40.75" resultid="7104" heatid="10496" lane="8" entrytime="00:00:41.33" entrycourse="LCM" />
                <RESULT eventid="1163" points="141" swimtime="00:03:53.85" resultid="7105" heatid="10553" lane="4" entrytime="00:03:43.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.35" />
                    <SPLIT distance="100" swimtime="00:01:43.89" />
                    <SPLIT distance="150" swimtime="00:02:49.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="241" swimtime="00:00:37.90" resultid="7106" heatid="10602" lane="5" entrytime="00:00:35.18" entrycourse="LCM" />
                <RESULT eventid="1297" points="201" swimtime="00:00:45.83" resultid="7107" heatid="10678" lane="0" entrytime="00:00:45.50" entrycourse="LCM" />
                <RESULT eventid="1333" points="145" swimtime="00:01:44.90" resultid="7108" heatid="10700" lane="9" entrytime="00:01:37.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Augusto Tafarel" birthdate="2009-12-23" gender="M" nation="BRA" license="423221" swrid="5820324" athleteid="7182" externalid="423221">
              <RESULTS>
                <RESULT eventid="1187" points="122" swimtime="00:00:52.30" resultid="7183" heatid="10570" lane="0" entrytime="00:00:52.27" entrycourse="LCM" />
                <RESULT eventid="1155" points="226" swimtime="00:01:16.17" resultid="7184" heatid="10539" lane="8" entrytime="00:01:16.25" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="De Reginalda" birthdate="2011-07-22" gender="M" nation="BRA" license="400323" swrid="5717257" athleteid="7138" externalid="400323">
              <RESULTS>
                <RESULT eventid="1103" points="396" swimtime="00:00:30.32" resultid="7139" heatid="10502" lane="1" />
                <RESULT eventid="1071" points="379" swimtime="00:02:34.53" resultid="7140" heatid="10477" lane="5" entrytime="00:02:36.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                    <SPLIT distance="100" swimtime="00:01:12.78" />
                    <SPLIT distance="150" swimtime="00:01:53.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="449" swimtime="00:01:00.58" resultid="7141" heatid="10547" lane="4" entrytime="00:01:01.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="469" swimtime="00:00:26.90" resultid="7142" heatid="10625" lane="0" entrytime="00:00:26.87" entrycourse="LCM" />
                <RESULT eventid="1305" points="430" swimtime="00:00:31.19" resultid="7143" heatid="10686" lane="0" entrytime="00:00:32.01" entrycourse="LCM" />
                <RESULT eventid="1373" points="416" swimtime="00:01:09.07" resultid="7144" heatid="10739" lane="1" entrytime="00:01:11.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Bernardi Iurk" birthdate="2012-04-14" gender="M" nation="BRA" license="408687" swrid="5725984" athleteid="7115" externalid="408687">
              <RESULTS>
                <RESULT eventid="1187" points="228" swimtime="00:00:42.43" resultid="7116" heatid="10570" lane="6" entrytime="00:00:46.63" entrycourse="LCM" />
                <RESULT eventid="1155" points="237" swimtime="00:01:14.96" resultid="7117" heatid="10539" lane="0" entrytime="00:01:16.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="239" swimtime="00:00:33.65" resultid="7118" heatid="10614" lane="5" entrytime="00:00:33.58" entrycourse="LCM" />
                <RESULT eventid="1219" points="211" swimtime="00:01:35.50" resultid="7119" heatid="10592" lane="6" entrytime="00:01:40.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="185" swimtime="00:02:58.81" resultid="7120" heatid="10661" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.78" />
                    <SPLIT distance="100" swimtime="00:01:22.63" />
                    <SPLIT distance="150" swimtime="00:02:10.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonia" lastname="Adam  Fracaro" birthdate="2010-04-27" gender="F" nation="BRA" license="382212" swrid="5588512" athleteid="7080" externalid="382212">
              <RESULTS>
                <RESULT eventid="1147" points="372" swimtime="00:01:11.88" resultid="7081" heatid="10528" lane="1" entrytime="00:01:13.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="390" swimtime="00:00:32.31" resultid="7082" heatid="10603" lane="7" entrytime="00:00:33.55" entrycourse="LCM" />
                <RESULT eventid="1281" points="337" swimtime="00:02:41.26" resultid="7083" heatid="10655" lane="1" entrytime="00:02:43.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.53" />
                    <SPLIT distance="100" swimtime="00:01:17.85" />
                    <SPLIT distance="150" swimtime="00:01:59.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="319" swimtime="00:05:44.31" resultid="7084" heatid="10713" lane="0" entrytime="00:05:47.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                    <SPLIT distance="100" swimtime="00:01:18.56" />
                    <SPLIT distance="150" swimtime="00:02:01.29" />
                    <SPLIT distance="200" swimtime="00:02:46.51" />
                    <SPLIT distance="250" swimtime="00:03:30.56" />
                    <SPLIT distance="300" swimtime="00:04:17.12" />
                    <SPLIT distance="350" swimtime="00:05:01.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="290" swimtime="00:01:26.26" resultid="7085" heatid="10728" lane="2" entrytime="00:01:27.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Zanchetta Silva" birthdate="2010-08-05" gender="F" nation="BRA" license="406865" swrid="5717308" athleteid="7151" externalid="406865">
              <RESULTS>
                <RESULT eventid="1147" points="245" swimtime="00:01:22.55" resultid="7152" heatid="10525" lane="5" entrytime="00:01:21.27" entrycourse="LCM" />
                <RESULT eventid="1227" status="DNS" swimtime="00:00:00.00" resultid="7153" heatid="10601" lane="4" entrytime="00:00:37.13" entrycourse="LCM" />
                <RESULT eventid="1297" points="216" swimtime="00:00:44.73" resultid="7154" heatid="10677" lane="4" entrytime="00:00:46.09" entrycourse="LCM" />
                <RESULT eventid="1365" points="183" swimtime="00:01:40.48" resultid="7155" heatid="10726" lane="5" entrytime="00:01:41.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabelly" lastname="Mendonca Bello" birthdate="2008-04-15" gender="F" nation="BRA" license="376996" swrid="5600217" athleteid="7093" externalid="376996" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1079" points="358" swimtime="00:03:13.54" resultid="7094" heatid="10484" lane="0" entrytime="00:03:07.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.14" />
                    <SPLIT distance="100" swimtime="00:01:29.97" />
                    <SPLIT distance="150" swimtime="00:02:20.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="446" swimtime="00:00:30.88" resultid="7095" heatid="10607" lane="3" entrytime="00:00:30.03" entrycourse="LCM" />
                <RESULT eventid="1211" points="366" swimtime="00:01:29.64" resultid="7096" heatid="10587" lane="4" entrytime="00:01:24.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="APAN-WS &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1323" points="264" swimtime="00:05:22.03" resultid="7187" heatid="10693" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                    <SPLIT distance="100" swimtime="00:01:16.83" />
                    <SPLIT distance="150" swimtime="00:02:00.26" />
                    <SPLIT distance="200" swimtime="00:02:53.14" />
                    <SPLIT distance="250" swimtime="00:03:29.20" />
                    <SPLIT distance="300" swimtime="00:04:11.49" />
                    <SPLIT distance="350" swimtime="00:04:43.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7170" number="1" />
                    <RELAYPOSITION athleteid="7115" number="2" />
                    <RELAYPOSITION athleteid="7145" number="3" />
                    <RELAYPOSITION athleteid="7109" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1391" points="301" swimtime="00:04:40.65" resultid="7188" heatid="10748" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                    <SPLIT distance="100" swimtime="00:01:05.85" />
                    <SPLIT distance="150" swimtime="00:01:40.38" />
                    <SPLIT distance="200" swimtime="00:02:20.42" />
                    <SPLIT distance="250" swimtime="00:02:52.63" />
                    <SPLIT distance="300" swimtime="00:03:29.90" />
                    <SPLIT distance="350" swimtime="00:04:02.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7145" number="1" />
                    <RELAYPOSITION athleteid="7115" number="2" />
                    <RELAYPOSITION athleteid="7170" number="3" />
                    <RELAYPOSITION athleteid="7109" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="F" name="APAN-WS &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1321" points="390" swimtime="00:05:14.04" resultid="7185" heatid="10692" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                    <SPLIT distance="100" swimtime="00:01:15.52" />
                    <SPLIT distance="150" swimtime="00:01:55.33" />
                    <SPLIT distance="200" swimtime="00:02:40.68" />
                    <SPLIT distance="250" swimtime="00:03:11.60" />
                    <SPLIT distance="300" swimtime="00:03:54.28" />
                    <SPLIT distance="350" swimtime="00:04:31.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7086" number="1" />
                    <RELAYPOSITION athleteid="7093" number="2" />
                    <RELAYPOSITION athleteid="7176" number="3" />
                    <RELAYPOSITION athleteid="7126" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1389" points="428" swimtime="00:04:35.87" resultid="7186" heatid="10747" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                    <SPLIT distance="100" swimtime="00:01:03.59" />
                    <SPLIT distance="150" swimtime="00:01:35.35" />
                    <SPLIT distance="200" swimtime="00:02:09.82" />
                    <SPLIT distance="250" swimtime="00:02:39.63" />
                    <SPLIT distance="300" swimtime="00:03:14.18" />
                    <SPLIT distance="350" swimtime="00:03:52.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7086" number="1" />
                    <RELAYPOSITION athleteid="7093" number="2" />
                    <RELAYPOSITION athleteid="7176" number="3" />
                    <RELAYPOSITION athleteid="7126" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="1007" nation="BRA" region="PR" clubid="9081" swrid="93785" name="Santa Mônica Clube De Campo" shortname="Santa Mônica">
          <ATHLETES>
            <ATHLETE firstname="Otto" lastname="Hedeke" birthdate="2011-03-24" gender="M" nation="BRA" license="372643" swrid="5588738" athleteid="9204" externalid="372643">
              <RESULTS>
                <RESULT eventid="1071" points="278" swimtime="00:02:51.30" resultid="9205" heatid="10474" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.64" />
                    <SPLIT distance="100" swimtime="00:01:21.29" />
                    <SPLIT distance="150" swimtime="00:02:06.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="395" swimtime="00:01:03.20" resultid="9206" heatid="10545" lane="1" entrytime="00:01:04.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="360" swimtime="00:00:29.37" resultid="9207" heatid="10615" lane="5" entrytime="00:00:32.43" entrycourse="LCM" />
                <RESULT eventid="1289" points="409" swimtime="00:02:17.36" resultid="9208" heatid="10669" lane="1" entrytime="00:02:20.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.27" />
                    <SPLIT distance="100" swimtime="00:01:06.12" />
                    <SPLIT distance="150" swimtime="00:01:42.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="402" swimtime="00:04:58.12" resultid="9209" heatid="10719" lane="4" entrytime="00:05:17.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.93" />
                    <SPLIT distance="100" swimtime="00:01:10.24" />
                    <SPLIT distance="150" swimtime="00:01:48.64" />
                    <SPLIT distance="200" swimtime="00:02:27.87" />
                    <SPLIT distance="250" swimtime="00:03:05.96" />
                    <SPLIT distance="300" swimtime="00:03:44.56" />
                    <SPLIT distance="350" swimtime="00:04:22.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Sofia Silva" birthdate="2007-05-28" gender="F" nation="BRA" license="390921" swrid="5600260" athleteid="9361" externalid="390921">
              <RESULTS>
                <RESULT eventid="1095" points="154" swimtime="00:00:45.51" resultid="9362" heatid="10495" lane="6" entrytime="00:00:45.47" entrycourse="LCM" />
                <RESULT eventid="1079" points="236" swimtime="00:03:42.31" resultid="9363" heatid="10482" lane="1" entrytime="00:03:42.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.39" />
                    <SPLIT distance="100" swimtime="00:01:44.16" />
                    <SPLIT distance="150" swimtime="00:02:43.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="251" swimtime="00:00:46.22" resultid="9364" heatid="10562" lane="7" entrytime="00:00:47.41" entrycourse="LCM" />
                <RESULT eventid="1211" points="257" swimtime="00:01:40.86" resultid="9365" heatid="10584" lane="0" entrytime="00:01:42.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="253" swimtime="00:00:42.46" resultid="9366" heatid="10677" lane="0" />
                <RESULT eventid="1265" points="253" swimtime="00:03:19.25" resultid="9367" heatid="10640" lane="8" entrytime="00:03:20.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.92" />
                    <SPLIT distance="100" swimtime="00:01:34.28" />
                    <SPLIT distance="150" swimtime="00:02:31.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emanuel" lastname="Correa Pertel Santos" birthdate="2010-09-15" gender="M" nation="BRA" license="421362" swrid="5810882" athleteid="9421" externalid="421362">
              <RESULTS>
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 11:13), Na chegada." eventid="1103" status="DSQ" swimtime="00:00:38.53" resultid="9422" heatid="10501" lane="0" />
                <RESULT eventid="1155" points="279" swimtime="00:01:11.00" resultid="9423" heatid="10541" lane="0" entrytime="00:01:12.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="258" swimtime="00:00:32.83" resultid="9424" heatid="10615" lane="1" entrytime="00:00:33.04" entrycourse="LCM" />
                <RESULT eventid="1289" points="268" swimtime="00:02:38.09" resultid="9425" heatid="10664" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                    <SPLIT distance="100" swimtime="00:01:12.24" />
                    <SPLIT distance="150" swimtime="00:01:54.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="De Siqueira Machado" birthdate="2012-05-25" gender="F" nation="BRA" license="377312" swrid="5588649" athleteid="9210" externalid="377312">
              <RESULTS>
                <RESULT comment="SW 10.2 - Não completou a distância total da prova.  (Horário: 10:01)" eventid="1079" status="DSQ" swimtime="00:00:00.00" resultid="9211" heatid="10481" lane="5" />
                <RESULT eventid="1179" points="362" swimtime="00:00:40.88" resultid="9212" heatid="10562" lane="6" entrytime="00:00:44.08" entrycourse="LCM" />
                <RESULT eventid="1147" points="296" swimtime="00:01:17.54" resultid="9213" heatid="10528" lane="0" entrytime="00:01:14.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="363" swimtime="00:00:33.08" resultid="9214" heatid="10604" lane="3" entrytime="00:00:31.96" entrycourse="LCM" />
                <RESULT eventid="1211" points="284" swimtime="00:01:37.52" resultid="9215" heatid="10584" lane="2" entrytime="00:01:38.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="301" swimtime="00:00:40.07" resultid="9216" heatid="10679" lane="3" entrytime="00:00:37.57" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Vianna" birthdate="2011-01-31" gender="M" nation="BRA" license="371380" swrid="5588947" athleteid="9197" externalid="371380">
              <RESULTS>
                <RESULT eventid="1123" points="403" swimtime="00:10:11.79" resultid="9198" heatid="10516" lane="4" entrytime="00:10:35.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                    <SPLIT distance="100" swimtime="00:01:13.51" />
                    <SPLIT distance="150" swimtime="00:01:52.25" />
                    <SPLIT distance="200" swimtime="00:02:30.53" />
                    <SPLIT distance="250" swimtime="00:03:08.76" />
                    <SPLIT distance="300" swimtime="00:03:48.24" />
                    <SPLIT distance="350" swimtime="00:04:27.19" />
                    <SPLIT distance="400" swimtime="00:05:07.36" />
                    <SPLIT distance="450" swimtime="00:05:46.58" />
                    <SPLIT distance="500" swimtime="00:06:25.94" />
                    <SPLIT distance="550" swimtime="00:07:04.59" />
                    <SPLIT distance="600" swimtime="00:07:44.52" />
                    <SPLIT distance="650" swimtime="00:08:22.35" />
                    <SPLIT distance="700" swimtime="00:09:00.13" />
                    <SPLIT distance="750" swimtime="00:09:35.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="333" swimtime="00:02:39.09" resultid="9199" heatid="10556" lane="2" entrytime="00:02:51.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                    <SPLIT distance="100" swimtime="00:01:14.20" />
                    <SPLIT distance="150" swimtime="00:01:57.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="404" swimtime="00:19:37.14" resultid="9200" heatid="10637" lane="4" entrytime="00:19:43.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                    <SPLIT distance="100" swimtime="00:01:13.82" />
                    <SPLIT distance="150" swimtime="00:01:51.85" />
                    <SPLIT distance="200" swimtime="00:02:31.84" />
                    <SPLIT distance="250" swimtime="00:03:09.52" />
                    <SPLIT distance="300" swimtime="00:03:49.72" />
                    <SPLIT distance="350" swimtime="00:04:28.27" />
                    <SPLIT distance="400" swimtime="00:05:08.22" />
                    <SPLIT distance="450" swimtime="00:05:46.84" />
                    <SPLIT distance="500" swimtime="00:06:27.31" />
                    <SPLIT distance="550" swimtime="00:07:07.08" />
                    <SPLIT distance="600" swimtime="00:07:47.87" />
                    <SPLIT distance="650" swimtime="00:08:26.25" />
                    <SPLIT distance="700" swimtime="00:09:06.86" />
                    <SPLIT distance="750" swimtime="00:09:46.62" />
                    <SPLIT distance="800" swimtime="00:10:26.57" />
                    <SPLIT distance="850" swimtime="00:11:05.29" />
                    <SPLIT distance="900" swimtime="00:11:46.47" />
                    <SPLIT distance="950" swimtime="00:12:25.96" />
                    <SPLIT distance="1000" swimtime="00:13:07.23" />
                    <SPLIT distance="1050" swimtime="00:13:47.20" />
                    <SPLIT distance="1100" swimtime="00:14:27.74" />
                    <SPLIT distance="1150" swimtime="00:15:07.12" />
                    <SPLIT distance="1200" swimtime="00:15:47.78" />
                    <SPLIT distance="1250" swimtime="00:16:26.70" />
                    <SPLIT distance="1300" swimtime="00:17:07.22" />
                    <SPLIT distance="1350" swimtime="00:17:45.22" />
                    <SPLIT distance="1400" swimtime="00:18:25.12" />
                    <SPLIT distance="1450" swimtime="00:19:00.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="406" swimtime="00:02:17.67" resultid="9201" heatid="10669" lane="0" entrytime="00:02:20.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                    <SPLIT distance="100" swimtime="00:01:06.57" />
                    <SPLIT distance="150" swimtime="00:01:42.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="363" swimtime="00:01:09.27" resultid="9202" heatid="10708" lane="1" entrytime="00:01:10.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="434" swimtime="00:04:50.62" resultid="9203" heatid="10720" lane="3" entrytime="00:05:00.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.73" />
                    <SPLIT distance="100" swimtime="00:01:09.78" />
                    <SPLIT distance="150" swimtime="00:01:47.45" />
                    <SPLIT distance="200" swimtime="00:02:25.42" />
                    <SPLIT distance="250" swimtime="00:03:01.61" />
                    <SPLIT distance="300" swimtime="00:03:38.70" />
                    <SPLIT distance="350" swimtime="00:04:15.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Marques" birthdate="2007-06-29" gender="M" nation="BRA" license="367257" swrid="5600213" athleteid="9312" externalid="367257">
              <RESULTS>
                <RESULT eventid="1123" points="345" swimtime="00:10:44.27" resultid="9313" heatid="10516" lane="5" entrytime="00:10:48.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="100" swimtime="00:01:12.07" />
                    <SPLIT distance="150" swimtime="00:01:50.71" />
                    <SPLIT distance="200" swimtime="00:02:30.40" />
                    <SPLIT distance="250" swimtime="00:03:09.35" />
                    <SPLIT distance="350" swimtime="00:04:29.41" />
                    <SPLIT distance="400" swimtime="00:05:09.48" />
                    <SPLIT distance="450" swimtime="00:05:51.50" />
                    <SPLIT distance="500" swimtime="00:06:32.35" />
                    <SPLIT distance="550" swimtime="00:07:14.83" />
                    <SPLIT distance="600" swimtime="00:07:54.70" />
                    <SPLIT distance="650" swimtime="00:08:37.82" />
                    <SPLIT distance="700" swimtime="00:09:20.67" />
                    <SPLIT distance="750" swimtime="00:10:01.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="331" swimtime="00:00:32.19" resultid="9314" heatid="10502" lane="8" />
                <RESULT eventid="1155" points="407" swimtime="00:01:02.58" resultid="9315" heatid="10546" lane="9" entrytime="00:01:03.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="397" swimtime="00:00:28.44" resultid="9316" heatid="10621" lane="8" entrytime="00:00:28.88" entrycourse="LCM" />
                <RESULT eventid="1289" points="393" swimtime="00:02:19.24" resultid="9317" heatid="10668" lane="4" entrytime="00:02:20.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                    <SPLIT distance="100" swimtime="00:01:07.36" />
                    <SPLIT distance="150" swimtime="00:01:43.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="380" swimtime="00:05:03.80" resultid="9318" heatid="10721" lane="9" entrytime="00:04:59.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                    <SPLIT distance="100" swimtime="00:01:10.90" />
                    <SPLIT distance="150" swimtime="00:01:49.00" />
                    <SPLIT distance="200" swimtime="00:02:28.31" />
                    <SPLIT distance="250" swimtime="00:03:07.02" />
                    <SPLIT distance="300" swimtime="00:03:46.92" />
                    <SPLIT distance="350" swimtime="00:04:26.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Marcos Morais" birthdate="2010-01-30" gender="M" nation="BRA" license="416736" swrid="5757093" athleteid="9334" externalid="416736">
              <RESULTS>
                <RESULT eventid="1071" points="289" swimtime="00:02:49.19" resultid="9335" heatid="10475" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.68" />
                    <SPLIT distance="100" swimtime="00:01:21.63" />
                    <SPLIT distance="150" swimtime="00:02:07.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="424" swimtime="00:00:34.54" resultid="9336" heatid="10573" lane="8" entrytime="00:00:36.39" entrycourse="LCM" />
                <RESULT eventid="1219" points="352" swimtime="00:01:20.53" resultid="9337" heatid="10597" lane="9" entrytime="00:01:18.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="326" swimtime="00:00:34.19" resultid="9338" heatid="10681" lane="7" />
                <RESULT eventid="1341" points="218" swimtime="00:01:22.13" resultid="9339" heatid="10703" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="324" swimtime="00:01:15.11" resultid="9340" heatid="10738" lane="1" entrytime="00:01:15.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caue" lastname="Sprengel Carneiro" birthdate="2004-07-12" gender="M" nation="BRA" license="324039" athleteid="9115" externalid="324039">
              <RESULTS>
                <RESULT eventid="1305" points="528" swimtime="00:00:29.12" resultid="9116" heatid="10682" lane="6" />
                <RESULT eventid="1373" points="506" swimtime="00:01:04.73" resultid="9117" heatid="10734" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Garay Costa" birthdate="2010-02-18" gender="M" nation="BRA" license="421361" swrid="5505752" athleteid="9415" externalid="421361">
              <RESULTS>
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 11:13), Na chegada." eventid="1103" status="DSQ" swimtime="00:00:37.94" resultid="9416" heatid="10501" lane="4" />
                <RESULT eventid="1155" points="327" swimtime="00:01:07.30" resultid="9417" heatid="10543" lane="1" entrytime="00:01:07.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="309" swimtime="00:00:30.90" resultid="9418" heatid="10618" lane="9" entrytime="00:00:30.92" entrycourse="LCM" />
                <RESULT eventid="1305" points="203" swimtime="00:00:40.02" resultid="9419" heatid="10683" lane="0" />
                <RESULT eventid="1289" points="311" swimtime="00:02:30.46" resultid="9420" heatid="10661" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.85" />
                    <SPLIT distance="100" swimtime="00:01:08.84" />
                    <SPLIT distance="150" swimtime="00:01:49.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Analyce" lastname="Nunes Porto Luz" birthdate="2006-10-29" gender="F" nation="BRA" license="369322" swrid="5600226" athleteid="9082" externalid="369322">
              <RESULTS>
                <RESULT eventid="1095" points="470" swimtime="00:00:31.41" resultid="9083" heatid="10498" lane="6" entrytime="00:00:31.37" entrycourse="LCM" />
                <RESULT eventid="1147" points="559" swimtime="00:01:02.75" resultid="9084" heatid="10534" lane="7" entrytime="00:01:03.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="512" swimtime="00:00:29.50" resultid="9085" heatid="10608" lane="5" entrytime="00:00:29.32" entrycourse="LCM" />
                <RESULT eventid="1297" points="454" swimtime="00:00:34.93" resultid="9086" heatid="10675" lane="4" />
                <RESULT eventid="1281" points="504" swimtime="00:02:20.98" resultid="9087" heatid="10660" lane="2" entrytime="00:02:18.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                    <SPLIT distance="100" swimtime="00:01:06.84" />
                    <SPLIT distance="150" swimtime="00:01:43.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="384" swimtime="00:01:15.89" resultid="9088" heatid="10702" lane="3" entrytime="00:01:11.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Pinterich Almeida" birthdate="2005-03-13" gender="M" nation="BRA" license="330749" swrid="5600235" athleteid="9118" externalid="330749">
              <RESULTS>
                <RESULT eventid="1235" points="584" swimtime="00:00:25.01" resultid="9119" heatid="10627" lane="7" entrytime="00:00:25.25" entrycourse="LCM" />
                <RESULT eventid="1305" points="516" swimtime="00:00:29.35" resultid="9120" heatid="10687" lane="6" entrytime="00:00:29.27" entrycourse="LCM" />
                <RESULT eventid="1289" points="545" swimtime="00:02:04.84" resultid="9121" heatid="10674" lane="5" entrytime="00:01:56.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.49" />
                    <SPLIT distance="100" swimtime="00:00:59.79" />
                    <SPLIT distance="150" swimtime="00:01:31.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="503" swimtime="00:01:02.17" resultid="9122" heatid="10711" lane="0" entrytime="00:01:00.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="509" swimtime="00:01:04.59" resultid="9123" heatid="10742" lane="2" entrytime="00:01:02.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="De Castro Paiva Maciel" birthdate="2008-04-10" gender="M" nation="BRA" license="378333" swrid="5622275" athleteid="9089" externalid="378333">
              <RESULTS>
                <RESULT eventid="1103" points="488" swimtime="00:00:28.27" resultid="9090" heatid="10507" lane="2" entrytime="00:00:28.33" entrycourse="LCM" />
                <RESULT eventid="1155" points="514" swimtime="00:00:57.91" resultid="9091" heatid="10549" lane="6" entrytime="00:00:58.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="456" swimtime="00:00:27.15" resultid="9092" heatid="10625" lane="9" entrytime="00:00:26.88" entrycourse="LCM" />
                <RESULT eventid="1305" points="368" swimtime="00:00:32.85" resultid="9093" heatid="10686" lane="8" entrytime="00:00:31.70" entrycourse="LCM" />
                <RESULT eventid="1289" points="495" swimtime="00:02:08.88" resultid="9094" heatid="10672" lane="5" entrytime="00:02:08.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.76" />
                    <SPLIT distance="100" swimtime="00:01:01.46" />
                    <SPLIT distance="150" swimtime="00:01:35.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="442" swimtime="00:01:04.91" resultid="9095" heatid="10709" lane="6" entrytime="00:01:05.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Larissa" lastname="Valera Mozzaquatro" birthdate="2012-10-13" gender="F" nation="BRA" license="421363" swrid="5810417" athleteid="9426" externalid="421363">
              <RESULTS>
                <RESULT eventid="1095" points="278" swimtime="00:00:37.39" resultid="9427" heatid="10494" lane="3" />
                <RESULT eventid="1063" points="357" swimtime="00:02:53.50" resultid="9428" heatid="10469" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="391" swimtime="00:01:10.71" resultid="9429" heatid="10529" lane="9" entrytime="00:01:12.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 9:42)" eventid="1227" status="DSQ" swimtime="00:00:32.26" resultid="9430" heatid="10605" lane="3" entrytime="00:00:31.28" entrycourse="LCM" />
                <RESULT eventid="1211" points="262" swimtime="00:01:40.14" resultid="9431" heatid="10584" lane="5" entrytime="00:01:37.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="353" swimtime="00:01:20.78" resultid="9432" heatid="10730" lane="9" entrytime="00:01:20.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Strapasson" birthdate="2012-03-01" gender="M" nation="BRA" license="371377" swrid="5602585" athleteid="9190" externalid="371377">
              <RESULTS>
                <RESULT eventid="1087" points="318" swimtime="00:03:03.82" resultid="9191" heatid="10489" lane="2" entrytime="00:03:06.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.91" />
                    <SPLIT distance="100" swimtime="00:01:27.11" />
                    <SPLIT distance="150" swimtime="00:02:15.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" status="WDR" swimtime="00:00:00.00" resultid="9192" />
                <RESULT eventid="1155" points="338" swimtime="00:01:06.61" resultid="9193" heatid="10544" lane="1" entrytime="00:01:06.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="372" swimtime="00:00:29.06" resultid="9194" heatid="10793" lane="4" entrytime="00:00:30.06" entrycourse="LCM" />
                <RESULT eventid="1219" points="299" swimtime="00:01:25.05" resultid="9195" heatid="10595" lane="7" entrytime="00:01:23.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="314" swimtime="00:02:29.91" resultid="9196" heatid="10666" lane="7" entrytime="00:02:36.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.80" />
                    <SPLIT distance="100" swimtime="00:01:11.34" />
                    <SPLIT distance="150" swimtime="00:01:51.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Augusto Vaz" birthdate="2011-06-25" gender="M" nation="BRA" license="401737" swrid="5661339" athleteid="9272" externalid="401737">
              <RESULTS>
                <RESULT eventid="1103" points="450" swimtime="00:00:29.05" resultid="9273" heatid="10506" lane="0" entrytime="00:00:30.92" entrycourse="LCM" />
                <RESULT eventid="1171" points="362" swimtime="00:02:34.73" resultid="9274" heatid="10557" lane="8" entrytime="00:02:36.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                    <SPLIT distance="100" swimtime="00:01:13.11" />
                    <SPLIT distance="150" swimtime="00:01:58.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="398" swimtime="00:00:28.41" resultid="9275" heatid="10622" lane="1" entrytime="00:00:28.22" entrycourse="LCM" />
                <RESULT eventid="1289" points="410" swimtime="00:02:17.27" resultid="9276" heatid="10668" lane="0" entrytime="00:02:25.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.11" />
                    <SPLIT distance="100" swimtime="00:01:05.85" />
                    <SPLIT distance="150" swimtime="00:01:42.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="473" swimtime="00:01:03.44" resultid="9277" heatid="10709" lane="5" entrytime="00:01:04.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="379" swimtime="00:05:04.07" resultid="9278" heatid="10718" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                    <SPLIT distance="100" swimtime="00:01:11.03" />
                    <SPLIT distance="150" swimtime="00:01:49.96" />
                    <SPLIT distance="200" swimtime="00:02:28.63" />
                    <SPLIT distance="250" swimtime="00:03:09.02" />
                    <SPLIT distance="300" swimtime="00:03:49.45" />
                    <SPLIT distance="350" swimtime="00:04:30.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edward" lastname="Luiz Santiago" birthdate="2012-02-02" gender="M" nation="BRA" license="413901" swrid="5742899" athleteid="9341" externalid="413901">
              <RESULTS>
                <RESULT eventid="1155" points="315" swimtime="00:01:08.18" resultid="9342" heatid="10542" lane="0" entrytime="00:01:10.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="311" swimtime="00:00:30.84" resultid="9343" heatid="10616" lane="1" entrytime="00:00:32.17" entrycourse="LCM" />
                <RESULT eventid="1305" points="242" swimtime="00:00:37.75" resultid="9344" heatid="10682" lane="4" />
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 16:27), Na volta dos 150m (Peito. Medley Individual)." eventid="1273" status="DSQ" swimtime="00:02:55.93" resultid="9345" heatid="10645" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.53" />
                    <SPLIT distance="100" swimtime="00:01:20.68" />
                    <SPLIT distance="150" swimtime="00:02:16.75" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 10.2 - Não completou a distância total da prova.  (Horário: 9:12)" eventid="1341" status="DSQ" swimtime="00:00:00.00" resultid="9346" heatid="10704" lane="1" />
                <RESULT eventid="1373" status="WDR" swimtime="00:00:00.00" resultid="9347" heatid="10736" lane="7" entrytime="00:01:21.96" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emily" lastname="Sayuri Tangueria De Lima" birthdate="2010-06-11" gender="F" nation="BRA" license="367215" swrid="5588901" athleteid="9180" externalid="367215">
              <RESULTS>
                <RESULT eventid="1095" points="412" swimtime="00:00:32.82" resultid="9181" heatid="10498" lane="8" entrytime="00:00:32.97" entrycourse="LCM" />
                <RESULT eventid="1163" points="334" swimtime="00:02:55.44" resultid="9182" heatid="10554" lane="2" entrytime="00:02:53.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.63" />
                    <SPLIT distance="100" swimtime="00:01:18.84" />
                    <SPLIT distance="150" swimtime="00:02:07.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="461" swimtime="00:01:06.89" resultid="9183" heatid="10531" lane="9" entrytime="00:01:07.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="452" swimtime="00:02:26.19" resultid="9184" heatid="10659" lane="1" entrytime="00:02:22.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                    <SPLIT distance="100" swimtime="00:01:10.63" />
                    <SPLIT distance="150" swimtime="00:01:49.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="412" swimtime="00:05:16.31" resultid="9185" heatid="10715" lane="3" entrytime="00:05:05.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                    <SPLIT distance="100" swimtime="00:01:15.21" />
                    <SPLIT distance="150" swimtime="00:01:55.44" />
                    <SPLIT distance="200" swimtime="00:02:36.29" />
                    <SPLIT distance="250" swimtime="00:03:16.02" />
                    <SPLIT distance="300" swimtime="00:03:56.60" />
                    <SPLIT distance="350" swimtime="00:04:38.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="391" swimtime="00:01:15.43" resultid="9186" heatid="10701" lane="4" entrytime="00:01:15.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietro" lastname="Lobo Mussoi" birthdate="2008-07-05" gender="M" nation="BRA" license="398573" swrid="5658061" athleteid="9395" externalid="398573">
              <RESULTS>
                <RESULT eventid="1123" points="366" swimtime="00:10:31.80" resultid="9396" heatid="10516" lane="6" entrytime="00:10:56.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                    <SPLIT distance="100" swimtime="00:01:09.69" />
                    <SPLIT distance="150" swimtime="00:01:48.26" />
                    <SPLIT distance="200" swimtime="00:02:27.62" />
                    <SPLIT distance="250" swimtime="00:03:07.40" />
                    <SPLIT distance="300" swimtime="00:03:47.69" />
                    <SPLIT distance="350" swimtime="00:04:28.26" />
                    <SPLIT distance="400" swimtime="00:05:10.00" />
                    <SPLIT distance="450" swimtime="00:05:50.27" />
                    <SPLIT distance="500" swimtime="00:06:32.17" />
                    <SPLIT distance="550" swimtime="00:07:13.66" />
                    <SPLIT distance="600" swimtime="00:07:53.91" />
                    <SPLIT distance="650" swimtime="00:08:34.07" />
                    <SPLIT distance="700" swimtime="00:09:13.90" />
                    <SPLIT distance="750" swimtime="00:09:52.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="498" swimtime="00:00:28.08" resultid="9397" heatid="10507" lane="9" entrytime="00:00:29.09" entrycourse="LCM" />
                <RESULT eventid="1155" points="491" swimtime="00:00:58.78" resultid="9398" heatid="10549" lane="9" entrytime="00:00:59.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="514" swimtime="00:00:26.10" resultid="9399" heatid="10626" lane="9" entrytime="00:00:26.09" entrycourse="LCM" />
                <RESULT eventid="1289" points="445" swimtime="00:02:13.55" resultid="9400" heatid="10663" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.47" />
                    <SPLIT distance="100" swimtime="00:01:01.62" />
                    <SPLIT distance="150" swimtime="00:01:37.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="440" swimtime="00:01:04.99" resultid="9401" heatid="10708" lane="5" entrytime="00:01:07.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Zattar" birthdate="2012-04-19" gender="F" nation="BRA" license="401736" swrid="5661351" athleteid="9265" externalid="401736">
              <RESULTS>
                <RESULT eventid="1079" points="363" swimtime="00:03:12.69" resultid="9266" heatid="10483" lane="6" entrytime="00:03:13.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.59" />
                    <SPLIT distance="100" swimtime="00:01:32.67" />
                    <SPLIT distance="150" swimtime="00:02:25.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="380" swimtime="00:00:40.23" resultid="9267" heatid="10563" lane="3" entrytime="00:00:40.80" entrycourse="LCM" />
                <RESULT eventid="1211" points="377" swimtime="00:01:28.70" resultid="9268" heatid="10585" lane="1" entrytime="00:01:32.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="380" swimtime="00:02:54.04" resultid="9269" heatid="10642" lane="0" entrytime="00:02:52.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                    <SPLIT distance="100" swimtime="00:01:20.48" />
                    <SPLIT distance="150" swimtime="00:02:15.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="411" swimtime="00:02:30.85" resultid="9270" heatid="10653" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                    <SPLIT distance="100" swimtime="00:01:12.64" />
                    <SPLIT distance="150" swimtime="00:01:52.61" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 8.2 - Braços não trazidos para frente simultaneamente sobre (em cima) a água.  (Horário: 8:59), SW 8.3 - Movimento alternado das pernas ou pés." eventid="1333" status="DSQ" swimtime="00:01:30.49" resultid="9271" heatid="10699" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Vitor Vicente" birthdate="2012-09-20" gender="M" nation="BRA" license="415246" swrid="5755345" athleteid="9328" externalid="415246">
              <RESULTS>
                <RESULT eventid="1087" points="176" swimtime="00:03:43.84" resultid="9329" heatid="10487" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.86" />
                    <SPLIT distance="100" swimtime="00:01:45.51" />
                    <SPLIT distance="150" swimtime="00:02:46.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="160" swimtime="00:00:47.71" resultid="9330" heatid="10570" lane="7" entrytime="00:00:48.23" entrycourse="LCM" />
                <RESULT eventid="1155" points="187" swimtime="00:01:21.02" resultid="9331" heatid="10538" lane="8" entrytime="00:01:24.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.4 - Movimentos das pernas não simultâneos.  (Horário: 9:24), Na volta dos 50m." eventid="1219" status="DSQ" swimtime="00:01:47.72" resultid="9332" heatid="10591" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="122" swimtime="00:00:47.41" resultid="9333" heatid="10683" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Larissa" lastname="Araujo Felix" birthdate="2010-05-27" gender="F" nation="BRA" license="393157" swrid="5622260" athleteid="9298" externalid="393157">
              <RESULTS>
                <RESULT eventid="1095" points="338" swimtime="00:00:35.05" resultid="9299" heatid="10496" lane="6" entrytime="00:00:37.19" entrycourse="LCM" />
                <RESULT eventid="1147" points="449" swimtime="00:01:07.52" resultid="9300" heatid="10530" lane="9" entrytime="00:01:09.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="431" swimtime="00:00:31.24" resultid="9301" heatid="10605" lane="7" entrytime="00:00:31.43" entrycourse="LCM" />
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 16:06), Na volta dos 150m (Peito. Medley Individual)." eventid="1265" status="DSQ" swimtime="00:03:03.17" resultid="9302" heatid="10640" lane="6" entrytime="00:03:13.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                    <SPLIT distance="100" swimtime="00:01:22.87" />
                    <SPLIT distance="150" swimtime="00:02:25.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="426" swimtime="00:02:29.13" resultid="9303" heatid="10657" lane="8" entrytime="00:02:29.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                    <SPLIT distance="100" swimtime="00:01:12.84" />
                    <SPLIT distance="150" swimtime="00:01:51.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="251" swimtime="00:01:27.45" resultid="9304" heatid="10700" lane="8" entrytime="00:01:31.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Araujo Farias" birthdate="2012-12-10" gender="F" nation="BRA" license="421354" swrid="5810904" athleteid="9409" externalid="421354">
              <RESULTS>
                <RESULT eventid="1179" points="142" swimtime="00:00:55.89" resultid="9410" heatid="10560" lane="5" />
                <RESULT eventid="1147" points="154" swimtime="00:01:36.44" resultid="9411" heatid="10524" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="183" swimtime="00:00:41.56" resultid="9412" heatid="10601" lane="7" entrytime="00:00:42.34" entrycourse="LCM" />
                <RESULT eventid="1211" points="153" swimtime="00:01:59.69" resultid="9413" heatid="10583" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="161" swimtime="00:03:26.03" resultid="9414" heatid="10654" lane="8" entrytime="00:03:25.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.77" />
                    <SPLIT distance="100" swimtime="00:01:42.29" />
                    <SPLIT distance="150" swimtime="00:02:35.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kauan" lastname="De Lima Dos Reis" birthdate="2010-04-18" gender="M" nation="BRA" license="413923" swrid="5811237" athleteid="9388" externalid="413923">
              <RESULTS>
                <RESULT eventid="1103" points="236" swimtime="00:00:36.00" resultid="9389" heatid="10500" lane="7" />
                <RESULT eventid="1087" points="246" swimtime="00:03:20.26" resultid="9390" heatid="10488" lane="5" entrytime="00:03:25.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.30" />
                    <SPLIT distance="100" swimtime="00:01:36.50" />
                    <SPLIT distance="150" swimtime="00:02:29.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="265" swimtime="00:00:40.36" resultid="9391" heatid="10567" lane="5" />
                <RESULT eventid="1155" points="286" swimtime="00:01:10.40" resultid="9392" heatid="10536" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="272" swimtime="00:00:32.26" resultid="9393" heatid="10616" lane="8" entrytime="00:00:32.19" entrycourse="LCM" />
                <RESULT eventid="1219" points="246" swimtime="00:01:30.69" resultid="9394" heatid="10593" lane="7" entrytime="00:01:32.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Larissa" lastname="Garcia Reschetti Rubbo" birthdate="2011-08-06" gender="F" nation="BRA" license="367053" swrid="5588720" athleteid="9131" externalid="367053" level="DCOMP IT">
              <RESULTS>
                <RESULT eventid="1079" points="356" swimtime="00:03:13.99" resultid="9132" heatid="10483" lane="7" entrytime="00:03:15.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.02" />
                    <SPLIT distance="100" swimtime="00:01:32.78" />
                    <SPLIT distance="150" swimtime="00:02:24.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="304" swimtime="00:00:43.32" resultid="9133" heatid="10562" lane="4" entrytime="00:00:43.09" entrycourse="LCM" />
                <RESULT eventid="1147" points="362" swimtime="00:01:12.52" resultid="9134" heatid="10528" lane="8" entrytime="00:01:14.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="350" swimtime="00:00:33.48" resultid="9135" heatid="10603" lane="6" entrytime="00:00:33.09" entrycourse="LCM" />
                <RESULT eventid="1211" points="324" swimtime="00:01:33.36" resultid="9136" heatid="10585" lane="5" entrytime="00:01:31.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="182" swimtime="00:01:37.23" resultid="9137" heatid="10700" lane="0" entrytime="00:01:35.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucca" lastname="Maceno Araujo" birthdate="2010-09-29" gender="M" nation="BRA" license="367056" swrid="5588788" athleteid="9145" externalid="367056">
              <RESULTS>
                <RESULT eventid="1103" points="450" swimtime="00:00:29.04" resultid="9146" heatid="10506" lane="4" entrytime="00:00:29.11" entrycourse="LCM" />
                <RESULT eventid="1171" points="317" swimtime="00:02:41.72" resultid="9147" heatid="10557" lane="0" entrytime="00:02:37.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                    <SPLIT distance="100" swimtime="00:01:12.90" />
                    <SPLIT distance="150" swimtime="00:01:56.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="419" swimtime="00:00:27.93" resultid="9148" heatid="10621" lane="6" entrytime="00:00:28.61" entrycourse="LCM" />
                <RESULT eventid="1289" points="431" swimtime="00:02:14.93" resultid="9149" heatid="10670" lane="8" entrytime="00:02:17.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                    <SPLIT distance="100" swimtime="00:01:04.44" />
                    <SPLIT distance="150" swimtime="00:01:39.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="442" swimtime="00:01:04.90" resultid="9150" heatid="10709" lane="2" entrytime="00:01:05.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="440" swimtime="00:04:49.28" resultid="9151" heatid="10722" lane="9" entrytime="00:04:50.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                    <SPLIT distance="100" swimtime="00:01:08.45" />
                    <SPLIT distance="150" swimtime="00:01:45.52" />
                    <SPLIT distance="200" swimtime="00:02:21.72" />
                    <SPLIT distance="250" swimtime="00:02:58.84" />
                    <SPLIT distance="300" swimtime="00:03:36.07" />
                    <SPLIT distance="350" swimtime="00:04:12.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathan" lastname="Torres Oliveira" birthdate="2008-04-10" gender="M" nation="BRA" license="400274" swrid="5653303" athleteid="9096" externalid="400274">
              <RESULTS>
                <RESULT eventid="1187" points="369" swimtime="00:00:36.16" resultid="9097" heatid="10572" lane="9" entrytime="00:00:39.96" entrycourse="LCM" />
                <RESULT eventid="1155" points="429" swimtime="00:01:01.49" resultid="9098" heatid="10548" lane="0" entrytime="00:01:00.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="469" swimtime="00:00:26.90" resultid="9099" heatid="10624" lane="7" entrytime="00:00:27.30" entrycourse="LCM" />
                <RESULT eventid="1289" points="389" swimtime="00:02:19.66" resultid="9100" heatid="10668" lane="7" entrytime="00:02:22.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                    <SPLIT distance="100" swimtime="00:01:07.92" />
                    <SPLIT distance="150" swimtime="00:01:45.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="342" swimtime="00:05:14.67" resultid="9101" heatid="10719" lane="3" entrytime="00:05:19.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                    <SPLIT distance="100" swimtime="00:01:10.91" />
                    <SPLIT distance="150" swimtime="00:01:51.65" />
                    <SPLIT distance="200" swimtime="00:02:34.17" />
                    <SPLIT distance="250" swimtime="00:03:16.80" />
                    <SPLIT distance="300" swimtime="00:03:59.84" />
                    <SPLIT distance="350" swimtime="00:04:38.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Nalle Bejes" birthdate="2010-04-20" gender="F" nation="BRA" license="377323" swrid="5588826" athleteid="9231" externalid="377323">
              <RESULTS>
                <RESULT eventid="1095" points="260" swimtime="00:00:38.26" resultid="9232" heatid="10495" lane="8" />
                <RESULT eventid="1079" points="391" swimtime="00:03:08.03" resultid="9233" heatid="10484" lane="2" entrytime="00:03:06.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.27" />
                    <SPLIT distance="100" swimtime="00:01:30.60" />
                    <SPLIT distance="150" swimtime="00:02:20.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="383" swimtime="00:00:40.15" resultid="9234" heatid="10563" lane="7" entrytime="00:00:41.50" entrycourse="LCM" />
                <RESULT eventid="1211" points="371" swimtime="00:01:29.23" resultid="9235" heatid="10587" lane="1" entrytime="00:01:25.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="399" swimtime="00:02:51.19" resultid="9236" heatid="10642" lane="2" entrytime="00:02:51.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.87" />
                    <SPLIT distance="100" swimtime="00:01:24.37" />
                    <SPLIT distance="150" swimtime="00:02:11.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="360" swimtime="00:05:30.80" resultid="9237" heatid="10714" lane="1" entrytime="00:05:23.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                    <SPLIT distance="100" swimtime="00:01:16.25" />
                    <SPLIT distance="150" swimtime="00:01:58.35" />
                    <SPLIT distance="200" swimtime="00:02:41.12" />
                    <SPLIT distance="250" swimtime="00:03:23.45" />
                    <SPLIT distance="300" swimtime="00:04:06.29" />
                    <SPLIT distance="350" swimtime="00:04:49.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Marques Machado" birthdate="2010-02-17" gender="M" nation="BRA" license="390918" swrid="5600212" athleteid="9245" externalid="390918">
              <RESULTS>
                <RESULT eventid="1123" points="430" swimtime="00:09:58.88" resultid="9246" heatid="10515" lane="6" entrytime="00:10:21.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.06" />
                    <SPLIT distance="100" swimtime="00:01:07.11" />
                    <SPLIT distance="150" swimtime="00:01:43.76" />
                    <SPLIT distance="200" swimtime="00:02:20.42" />
                    <SPLIT distance="250" swimtime="00:02:57.11" />
                    <SPLIT distance="300" swimtime="00:03:35.52" />
                    <SPLIT distance="350" swimtime="00:04:13.57" />
                    <SPLIT distance="400" swimtime="00:04:51.95" />
                    <SPLIT distance="450" swimtime="00:05:31.30" />
                    <SPLIT distance="500" swimtime="00:06:10.67" />
                    <SPLIT distance="550" swimtime="00:06:49.00" />
                    <SPLIT distance="600" swimtime="00:07:28.09" />
                    <SPLIT distance="650" swimtime="00:08:07.55" />
                    <SPLIT distance="700" swimtime="00:08:46.27" />
                    <SPLIT distance="750" swimtime="00:09:23.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="371" swimtime="00:00:30.99" resultid="9247" heatid="10505" lane="4" entrytime="00:00:31.06" entrycourse="LCM" />
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 19:02), 150m" eventid="1171" status="DSQ" swimtime="00:02:42.85" resultid="9248" heatid="10557" lane="9" entrytime="00:02:40.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                    <SPLIT distance="100" swimtime="00:01:16.21" />
                    <SPLIT distance="150" swimtime="00:02:00.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="423" swimtime="00:19:19.31" resultid="9249" heatid="10636" lane="2" entrytime="00:19:09.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="100" swimtime="00:01:09.47" />
                    <SPLIT distance="150" swimtime="00:01:47.12" />
                    <SPLIT distance="200" swimtime="00:02:25.72" />
                    <SPLIT distance="250" swimtime="00:03:04.46" />
                    <SPLIT distance="300" swimtime="00:03:43.01" />
                    <SPLIT distance="350" swimtime="00:04:20.83" />
                    <SPLIT distance="400" swimtime="00:04:59.96" />
                    <SPLIT distance="450" swimtime="00:05:38.54" />
                    <SPLIT distance="500" swimtime="00:06:18.61" />
                    <SPLIT distance="550" swimtime="00:06:57.57" />
                    <SPLIT distance="600" swimtime="00:07:36.06" />
                    <SPLIT distance="650" swimtime="00:08:14.70" />
                    <SPLIT distance="700" swimtime="00:08:53.49" />
                    <SPLIT distance="750" swimtime="00:09:32.28" />
                    <SPLIT distance="800" swimtime="00:10:11.64" />
                    <SPLIT distance="850" swimtime="00:10:50.82" />
                    <SPLIT distance="900" swimtime="00:11:30.40" />
                    <SPLIT distance="950" swimtime="00:12:09.66" />
                    <SPLIT distance="1000" swimtime="00:12:49.57" />
                    <SPLIT distance="1050" swimtime="00:13:29.10" />
                    <SPLIT distance="1100" swimtime="00:14:08.57" />
                    <SPLIT distance="1150" swimtime="00:14:47.86" />
                    <SPLIT distance="1200" swimtime="00:15:28.11" />
                    <SPLIT distance="1250" swimtime="00:16:07.61" />
                    <SPLIT distance="1300" swimtime="00:16:46.96" />
                    <SPLIT distance="1350" swimtime="00:17:25.52" />
                    <SPLIT distance="1400" swimtime="00:18:05.14" />
                    <SPLIT distance="1450" swimtime="00:18:44.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="426" swimtime="00:02:15.47" resultid="9250" heatid="10669" lane="2" entrytime="00:02:19.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                    <SPLIT distance="100" swimtime="00:01:05.47" />
                    <SPLIT distance="150" swimtime="00:01:41.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="400" swimtime="00:04:58.44" resultid="9251" heatid="10720" lane="5" entrytime="00:04:59.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                    <SPLIT distance="100" swimtime="00:01:07.95" />
                    <SPLIT distance="150" swimtime="00:01:44.96" />
                    <SPLIT distance="200" swimtime="00:02:23.33" />
                    <SPLIT distance="250" swimtime="00:03:01.66" />
                    <SPLIT distance="300" swimtime="00:03:40.40" />
                    <SPLIT distance="350" swimtime="00:04:19.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Murara" birthdate="1991-04-12" gender="M" nation="BRA" license="386866" swrid="5622296" athleteid="9319" externalid="386866">
              <RESULTS>
                <RESULT eventid="1235" points="548" swimtime="00:00:25.54" resultid="9320" heatid="10627" lane="5" entrytime="00:00:25.12" entrycourse="LCM" />
                <RESULT eventid="1305" points="517" swimtime="00:00:29.32" resultid="9321" heatid="10687" lane="4" entrytime="00:00:28.58" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luan" lastname="Felipe Ribeiro" birthdate="2010-11-05" gender="M" nation="BRA" license="423888" swrid="5820333" athleteid="9455" externalid="423888">
              <RESULTS>
                <RESULT eventid="1103" points="283" swimtime="00:00:33.90" resultid="9456" heatid="10500" lane="2" />
                <RESULT eventid="1187" points="285" swimtime="00:00:39.41" resultid="9457" heatid="10567" lane="2" />
                <RESULT eventid="1155" points="342" swimtime="00:01:06.34" resultid="9458" heatid="10537" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="337" swimtime="00:00:30.03" resultid="9459" heatid="10610" lane="3" />
                <RESULT eventid="1289" points="307" swimtime="00:02:31.10" resultid="9460" heatid="10664" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                    <SPLIT distance="100" swimtime="00:01:10.38" />
                    <SPLIT distance="150" swimtime="00:01:50.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="271" swimtime="00:05:39.89" resultid="9461" heatid="10718" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.77" />
                    <SPLIT distance="100" swimtime="00:01:16.58" />
                    <SPLIT distance="150" swimtime="00:01:59.52" />
                    <SPLIT distance="200" swimtime="00:02:43.88" />
                    <SPLIT distance="250" swimtime="00:03:28.12" />
                    <SPLIT distance="300" swimtime="00:04:13.23" />
                    <SPLIT distance="350" swimtime="00:04:56.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Gabriel Camargo" birthdate="2010-07-03" gender="M" nation="BRA" license="421421" swrid="4199554" athleteid="9442" externalid="421421">
              <RESULTS>
                <RESULT eventid="1103" points="254" swimtime="00:00:35.12" resultid="9443" heatid="10501" lane="3" />
                <RESULT eventid="1155" points="310" swimtime="00:01:08.50" resultid="9444" heatid="10542" lane="5" entrytime="00:01:08.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="286" swimtime="00:00:31.72" resultid="9445" heatid="10616" lane="2" entrytime="00:00:32.02" entrycourse="LCM" />
                <RESULT eventid="1289" points="295" swimtime="00:02:33.09" resultid="9446" heatid="10667" lane="0" entrytime="00:02:30.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                    <SPLIT distance="100" swimtime="00:01:13.29" />
                    <SPLIT distance="150" swimtime="00:01:54.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="298" swimtime="00:05:29.20" resultid="9447" heatid="10718" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                    <SPLIT distance="100" swimtime="00:01:17.19" />
                    <SPLIT distance="150" swimtime="00:01:59.91" />
                    <SPLIT distance="200" swimtime="00:02:42.11" />
                    <SPLIT distance="250" swimtime="00:03:25.66" />
                    <SPLIT distance="300" swimtime="00:04:08.85" />
                    <SPLIT distance="350" swimtime="00:04:50.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carol" lastname="Nalle Bejes" birthdate="2010-04-20" gender="F" nation="BRA" license="377315" swrid="5588824" athleteid="9217" externalid="377315">
              <RESULTS>
                <RESULT eventid="1079" points="459" swimtime="00:02:58.24" resultid="9218" heatid="10486" lane="0" entrytime="00:02:56.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.67" />
                    <SPLIT distance="100" swimtime="00:01:25.89" />
                    <SPLIT distance="150" swimtime="00:02:13.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="434" swimtime="00:00:38.50" resultid="9219" heatid="10565" lane="8" entrytime="00:00:37.14" entrycourse="LCM" />
                <RESULT eventid="1211" points="452" swimtime="00:01:23.56" resultid="9220" heatid="10588" lane="0" entrytime="00:01:23.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="383" swimtime="00:02:53.52" resultid="9221" heatid="10639" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.29" />
                    <SPLIT distance="100" swimtime="00:01:27.22" />
                    <SPLIT distance="150" swimtime="00:02:14.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="445" swimtime="00:02:27.00" resultid="9222" heatid="10658" lane="1" entrytime="00:02:26.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                    <SPLIT distance="100" swimtime="00:01:11.09" />
                    <SPLIT distance="150" swimtime="00:01:49.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="401" swimtime="00:05:19.04" resultid="9223" heatid="10714" lane="5" entrytime="00:05:14.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                    <SPLIT distance="100" swimtime="00:01:12.47" />
                    <SPLIT distance="150" swimtime="00:01:51.81" />
                    <SPLIT distance="200" swimtime="00:02:32.34" />
                    <SPLIT distance="250" swimtime="00:03:13.93" />
                    <SPLIT distance="300" swimtime="00:03:57.56" />
                    <SPLIT distance="350" swimtime="00:04:40.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Mosko Oliveira" birthdate="2009-01-07" gender="M" nation="BRA" license="421418" swrid="5820328" athleteid="9438" externalid="421418">
              <RESULTS>
                <RESULT eventid="1155" points="417" swimtime="00:01:02.10" resultid="9439" heatid="10537" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="401" swimtime="00:00:28.34" resultid="9440" heatid="10621" lane="0" entrytime="00:00:28.94" entrycourse="LCM" />
                <RESULT eventid="1289" points="357" swimtime="00:02:23.73" resultid="9441" heatid="10662" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                    <SPLIT distance="100" swimtime="00:01:06.62" />
                    <SPLIT distance="150" swimtime="00:01:45.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Cavassin Ieger" birthdate="2011-08-31" gender="M" nation="BRA" license="367149" swrid="5588743" athleteid="9159" externalid="367149">
              <RESULTS>
                <RESULT eventid="1103" points="326" swimtime="00:00:32.35" resultid="9160" heatid="10500" lane="1" />
                <RESULT eventid="1087" points="354" swimtime="00:02:57.29" resultid="9161" heatid="10490" lane="0" entrytime="00:02:58.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                    <SPLIT distance="100" swimtime="00:01:23.82" />
                    <SPLIT distance="150" swimtime="00:02:09.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="379" swimtime="00:00:35.84" resultid="9162" heatid="10573" lane="7" entrytime="00:00:36.09" entrycourse="LCM" />
                <RESULT eventid="1235" points="335" swimtime="00:00:30.08" resultid="9163" heatid="10611" lane="9" />
                <RESULT eventid="1219" points="370" swimtime="00:01:19.17" resultid="9164" heatid="10596" lane="2" entrytime="00:01:19.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="339" swimtime="00:02:43.43" resultid="9165" heatid="10649" lane="0" entrytime="00:02:43.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="100" swimtime="00:01:19.77" />
                    <SPLIT distance="150" swimtime="00:02:04.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luisa" lastname="Hoch Santos" birthdate="2011-07-05" gender="F" nation="BRA" license="403784" swrid="5684570" athleteid="9286" externalid="403784">
              <RESULTS>
                <RESULT eventid="1095" points="110" swimtime="00:00:50.95" resultid="9287" heatid="10495" lane="0" />
                <RESULT eventid="1147" points="242" swimtime="00:01:22.94" resultid="9288" heatid="10525" lane="7" entrytime="00:01:25.21" entrycourse="LCM" />
                <RESULT eventid="1227" points="265" swimtime="00:00:36.74" resultid="9289" heatid="10601" lane="6" entrytime="00:00:38.20" entrycourse="LCM" />
                <RESULT eventid="1297" points="211" swimtime="00:00:45.09" resultid="9290" heatid="10677" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Bello Costa Lange" birthdate="2010-09-13" gender="M" nation="BRA" license="367152" swrid="5588547" athleteid="9173" externalid="367152">
              <RESULTS>
                <RESULT eventid="1103" points="407" swimtime="00:00:30.04" resultid="9174" heatid="10505" lane="1" entrytime="00:00:31.96" entrycourse="LCM" />
                <RESULT eventid="1087" points="427" swimtime="00:02:46.61" resultid="9175" heatid="10491" lane="1" entrytime="00:02:48.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.78" />
                    <SPLIT distance="100" swimtime="00:01:18.35" />
                    <SPLIT distance="150" swimtime="00:02:03.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="437" swimtime="00:00:34.19" resultid="9176" heatid="10574" lane="8" entrytime="00:00:35.02" entrycourse="LCM" />
                <RESULT eventid="1219" points="443" swimtime="00:01:14.57" resultid="9177" heatid="10597" lane="2" entrytime="00:01:15.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 8.3 - Movimento alternado das pernas ou pés.  (Horário: 16:51), Durante o percurso (Borboleta, Medley Individual)." eventid="1273" status="DSQ" swimtime="00:02:31.11" resultid="9178" heatid="10650" lane="0" entrytime="00:02:34.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                    <SPLIT distance="100" swimtime="00:01:14.23" />
                    <SPLIT distance="150" swimtime="00:01:55.62" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 8.3 - Movimento alternado das pernas ou pés.  (Horário: 9:19)" eventid="1341" status="DSQ" swimtime="00:01:10.32" resultid="9179" heatid="10707" lane="1" entrytime="00:01:13.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexandre" lastname="Celli Schneider" birthdate="2011-02-21" gender="M" nation="BRA" license="367055" swrid="5588587" athleteid="9138" externalid="367055">
              <RESULTS>
                <RESULT eventid="1071" points="419" swimtime="00:02:29.49" resultid="9139" heatid="10478" lane="0" entrytime="00:02:33.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                    <SPLIT distance="100" swimtime="00:01:13.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="372" swimtime="00:02:33.40" resultid="9140" heatid="10557" lane="7" entrytime="00:02:36.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.51" />
                    <SPLIT distance="100" swimtime="00:01:14.12" />
                    <SPLIT distance="150" swimtime="00:01:55.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="440" swimtime="00:00:30.96" resultid="9141" heatid="10685" lane="4" entrytime="00:00:32.59" entrycourse="LCM" />
                <RESULT eventid="1273" points="438" swimtime="00:02:30.02" resultid="9142" heatid="10649" lane="7" entrytime="00:02:42.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                    <SPLIT distance="100" swimtime="00:01:10.97" />
                    <SPLIT distance="150" swimtime="00:01:56.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="410" swimtime="00:01:06.56" resultid="9143" heatid="10709" lane="0" entrytime="00:01:07.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="459" swimtime="00:01:06.87" resultid="9144" heatid="10739" lane="2" entrytime="00:01:10.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Freitas Szucs" birthdate="2011-10-02" gender="M" nation="BRA" license="377272" swrid="5588708" athleteid="9374" externalid="377272">
              <RESULTS>
                <RESULT eventid="1103" points="237" swimtime="00:00:35.98" resultid="9375" heatid="10503" lane="1" entrytime="00:00:36.67" entrycourse="LCM" />
                <RESULT eventid="1187" points="191" swimtime="00:00:45.02" resultid="9376" heatid="10569" lane="9" />
                <RESULT eventid="1155" points="271" swimtime="00:01:11.69" resultid="9377" heatid="10541" lane="2" entrytime="00:01:11.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="282" swimtime="00:00:31.88" resultid="9378" heatid="10615" lane="6" entrytime="00:00:32.52" entrycourse="LCM" />
                <RESULT eventid="1305" points="145" swimtime="00:00:44.76" resultid="9379" heatid="10682" lane="5" />
                <RESULT eventid="1289" points="243" swimtime="00:02:43.40" resultid="9380" heatid="10665" lane="0" entrytime="00:02:50.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                    <SPLIT distance="100" swimtime="00:01:18.81" />
                    <SPLIT distance="150" swimtime="00:02:02.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natália" lastname="Bacellar" birthdate="2011-02-01" gender="F" nation="BRA" license="386865" swrid="5810964" athleteid="9355" externalid="386865">
              <RESULTS>
                <RESULT eventid="1179" points="188" swimtime="00:00:50.88" resultid="9356" heatid="10561" lane="4" entrytime="00:00:53.63" entrycourse="LCM" />
                <RESULT eventid="1147" points="192" swimtime="00:01:29.49" resultid="9357" heatid="10525" lane="1" entrytime="00:01:34.18" entrycourse="LCM" />
                <RESULT eventid="1227" points="165" swimtime="00:00:42.96" resultid="9358" heatid="10601" lane="2" entrytime="00:00:40.15" entrycourse="LCM" />
                <RESULT eventid="1211" points="160" swimtime="00:01:58.02" resultid="9359" heatid="10583" lane="5" entrytime="00:01:52.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="180" swimtime="00:00:47.50" resultid="9360" heatid="10676" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Luiz Cruz" birthdate="2012-10-13" gender="M" nation="BRA" license="393209" swrid="5616447" athleteid="9252" externalid="393209">
              <RESULTS>
                <RESULT eventid="1155" points="220" swimtime="00:01:16.80" resultid="9253" heatid="10538" lane="4" entrytime="00:01:19.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="217" swimtime="00:00:34.75" resultid="9254" heatid="10614" lane="7" entrytime="00:00:34.91" entrycourse="LCM" />
                <RESULT eventid="1219" points="140" swimtime="00:01:49.36" resultid="9255" heatid="10592" lane="0" entrytime="00:01:43.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="210" swimtime="00:02:51.37" resultid="9256" heatid="10664" lane="4" entrytime="00:02:54.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.82" />
                    <SPLIT distance="100" swimtime="00:01:19.87" />
                    <SPLIT distance="150" swimtime="00:02:06.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="112" swimtime="00:01:42.58" resultid="9257" heatid="10704" lane="5" entrytime="00:01:50.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Blansky Hagebock" birthdate="2008-08-15" gender="M" nation="BRA" license="339123" swrid="5455418" athleteid="9109" externalid="339123">
              <RESULTS>
                <RESULT eventid="1103" points="496" swimtime="00:00:28.13" resultid="9110" heatid="10507" lane="8" entrytime="00:00:28.79" entrycourse="LCM" />
                <RESULT eventid="1155" points="570" swimtime="00:00:55.95" resultid="9111" heatid="10551" lane="7" entrytime="00:00:55.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="534" swimtime="00:00:25.77" resultid="9112" heatid="10626" lane="6" entrytime="00:00:25.73" entrycourse="LCM" />
                <RESULT eventid="1289" points="487" swimtime="00:02:09.59" resultid="9113" heatid="10672" lane="7" entrytime="00:02:09.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.40" />
                    <SPLIT distance="100" swimtime="00:01:02.61" />
                    <SPLIT distance="150" swimtime="00:01:37.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="462" swimtime="00:04:44.49" resultid="9114" heatid="10722" lane="5" entrytime="00:04:42.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                    <SPLIT distance="100" swimtime="00:01:06.33" />
                    <SPLIT distance="150" swimtime="00:01:42.25" />
                    <SPLIT distance="200" swimtime="00:02:18.53" />
                    <SPLIT distance="250" swimtime="00:02:55.06" />
                    <SPLIT distance="300" swimtime="00:03:32.24" />
                    <SPLIT distance="350" swimtime="00:04:09.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Goncalves Plocharski" birthdate="2011-08-01" gender="M" nation="BRA" license="413922" swrid="5811244" athleteid="9348" externalid="413922">
              <RESULTS>
                <RESULT eventid="1087" points="244" swimtime="00:03:20.63" resultid="9349" heatid="10487" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.17" />
                    <SPLIT distance="100" swimtime="00:01:35.70" />
                    <SPLIT distance="150" swimtime="00:02:30.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="260" swimtime="00:00:40.65" resultid="9350" heatid="10569" lane="7" />
                <RESULT eventid="1155" points="240" swimtime="00:01:14.59" resultid="9351" heatid="10536" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="268" swimtime="00:01:28.18" resultid="9352" heatid="10591" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="207" swimtime="00:00:39.75" resultid="9353" heatid="10684" lane="2" entrytime="00:00:38.55" entrycourse="LCM" />
                <RESULT eventid="1373" points="198" swimtime="00:01:28.44" resultid="9354" heatid="10734" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Diego" lastname="Brasil Caropreso" birthdate="2009-10-29" gender="M" nation="BRA" license="399502" swrid="5653287" athleteid="9291" externalid="399502">
              <RESULTS>
                <RESULT eventid="1103" points="389" swimtime="00:00:30.49" resultid="9292" heatid="10505" lane="2" entrytime="00:00:31.69" entrycourse="LCM" />
                <RESULT eventid="1155" points="466" swimtime="00:00:59.81" resultid="9293" heatid="10548" lane="1" entrytime="00:01:00.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="416" swimtime="00:00:28.01" resultid="9294" heatid="10623" lane="0" entrytime="00:00:27.80" entrycourse="LCM" />
                <RESULT eventid="1289" points="408" swimtime="00:02:17.42" resultid="9295" heatid="10670" lane="2" entrytime="00:02:16.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                    <SPLIT distance="100" swimtime="00:01:03.97" />
                    <SPLIT distance="150" swimtime="00:01:40.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="297" swimtime="00:01:14.08" resultid="9296" heatid="10706" lane="2" entrytime="00:01:17.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="384" swimtime="00:05:02.54" resultid="9297" heatid="10721" lane="8" entrytime="00:04:58.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                    <SPLIT distance="100" swimtime="00:01:11.28" />
                    <SPLIT distance="150" swimtime="00:01:50.87" />
                    <SPLIT distance="200" swimtime="00:02:29.65" />
                    <SPLIT distance="250" swimtime="00:03:09.11" />
                    <SPLIT distance="300" swimtime="00:03:46.72" />
                    <SPLIT distance="350" swimtime="00:04:28.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathan" lastname="Cordeiro Pimentel" birthdate="2012-04-30" gender="M" nation="BRA" license="421364" swrid="5806843" athleteid="9433" externalid="421364">
              <RESULTS>
                <RESULT eventid="1187" points="165" swimtime="00:00:47.30" resultid="9434" heatid="10567" lane="8" />
                <RESULT eventid="1155" points="183" swimtime="00:01:21.68" resultid="9435" heatid="10538" lane="7" entrytime="00:01:22.98" entrycourse="LCM" />
                <RESULT eventid="1235" points="195" swimtime="00:00:36.05" resultid="9436" heatid="10614" lane="1" entrytime="00:00:35.36" entrycourse="LCM" />
                <RESULT eventid="1305" points="152" swimtime="00:00:44.09" resultid="9437" heatid="10681" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Wenceslau Bitencourt" birthdate="2012-02-11" gender="M" nation="BRA" license="377318" swrid="5602591" athleteid="9224" externalid="377318">
              <RESULTS>
                <RESULT eventid="1103" status="WDR" swimtime="00:00:00.00" resultid="9225" heatid="10503" lane="7" entrytime="00:00:36.14" entrycourse="LCM" />
                <RESULT eventid="1155" status="WDR" swimtime="00:00:00.00" resultid="9226" heatid="10539" lane="6" entrytime="00:01:14.86" entrycourse="LCM" />
                <RESULT eventid="1235" status="WDR" swimtime="00:00:00.00" resultid="9227" heatid="10615" lane="7" entrytime="00:00:32.66" entrycourse="LCM" />
                <RESULT eventid="1273" status="WDR" swimtime="00:00:00.00" resultid="9228" heatid="10647" lane="6" entrytime="00:02:56.42" entrycourse="LCM" />
                <RESULT eventid="1289" status="WDR" swimtime="00:00:00.00" resultid="9229" heatid="10666" lane="4" entrytime="00:02:33.82" entrycourse="LCM" />
                <RESULT eventid="1341" status="WDR" swimtime="00:00:00.00" resultid="9230" heatid="10706" lane="1" entrytime="00:01:18.31" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Victor Dallastra" birthdate="2010-08-21" gender="M" nation="BRA" license="408024" swrid="5723028" athleteid="9322" externalid="408024">
              <RESULTS>
                <RESULT eventid="1103" points="404" swimtime="00:00:30.11" resultid="9323" heatid="10505" lane="8" entrytime="00:00:32.04" entrycourse="LCM" />
                <RESULT eventid="1155" points="491" swimtime="00:00:58.79" resultid="9324" heatid="10549" lane="2" entrytime="00:00:58.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="427" swimtime="00:00:27.76" resultid="9325" heatid="10624" lane="0" entrytime="00:00:27.40" entrycourse="LCM" />
                <RESULT eventid="1289" points="512" swimtime="00:02:07.50" resultid="9326" heatid="10672" lane="2" entrytime="00:02:09.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.94" />
                    <SPLIT distance="100" swimtime="00:01:01.55" />
                    <SPLIT distance="150" swimtime="00:01:35.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="518" swimtime="00:04:33.94" resultid="9327" heatid="10723" lane="6" entrytime="00:04:33.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.77" />
                    <SPLIT distance="100" swimtime="00:01:03.40" />
                    <SPLIT distance="150" swimtime="00:01:38.00" />
                    <SPLIT distance="200" swimtime="00:02:13.35" />
                    <SPLIT distance="250" swimtime="00:02:48.96" />
                    <SPLIT distance="300" swimtime="00:03:25.34" />
                    <SPLIT distance="350" swimtime="00:04:01.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kedny" lastname="Correa" birthdate="2004-11-05" gender="M" nation="BRA" license="383858" swrid="5600142" athleteid="9381" externalid="383858">
              <RESULTS>
                <RESULT eventid="1123" points="440" swimtime="00:09:54.36" resultid="9382" heatid="10514" lane="1" entrytime="00:09:54.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.66" />
                    <SPLIT distance="100" swimtime="00:01:08.05" />
                    <SPLIT distance="150" swimtime="00:01:43.83" />
                    <SPLIT distance="200" swimtime="00:02:20.63" />
                    <SPLIT distance="250" swimtime="00:02:57.19" />
                    <SPLIT distance="300" swimtime="00:03:34.59" />
                    <SPLIT distance="350" swimtime="00:04:11.86" />
                    <SPLIT distance="400" swimtime="00:04:49.78" />
                    <SPLIT distance="450" swimtime="00:05:27.50" />
                    <SPLIT distance="500" swimtime="00:06:05.71" />
                    <SPLIT distance="550" swimtime="00:06:44.07" />
                    <SPLIT distance="600" swimtime="00:07:22.70" />
                    <SPLIT distance="650" swimtime="00:08:00.61" />
                    <SPLIT distance="700" swimtime="00:08:39.29" />
                    <SPLIT distance="750" swimtime="00:09:16.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="282" swimtime="00:02:48.26" resultid="9383" heatid="10556" lane="6" entrytime="00:02:46.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                    <SPLIT distance="100" swimtime="00:01:12.01" />
                    <SPLIT distance="150" swimtime="00:01:57.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="472" swimtime="00:18:37.70" resultid="9384" heatid="10636" lane="4" entrytime="00:18:36.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                    <SPLIT distance="100" swimtime="00:01:08.65" />
                    <SPLIT distance="150" swimtime="00:01:45.36" />
                    <SPLIT distance="200" swimtime="00:02:22.55" />
                    <SPLIT distance="250" swimtime="00:02:59.93" />
                    <SPLIT distance="300" swimtime="00:03:37.74" />
                    <SPLIT distance="350" swimtime="00:04:15.10" />
                    <SPLIT distance="400" swimtime="00:04:52.84" />
                    <SPLIT distance="450" swimtime="00:05:30.44" />
                    <SPLIT distance="500" swimtime="00:06:08.68" />
                    <SPLIT distance="550" swimtime="00:06:45.62" />
                    <SPLIT distance="600" swimtime="00:07:23.23" />
                    <SPLIT distance="650" swimtime="00:08:00.20" />
                    <SPLIT distance="700" swimtime="00:08:37.76" />
                    <SPLIT distance="750" swimtime="00:09:14.50" />
                    <SPLIT distance="800" swimtime="00:09:52.14" />
                    <SPLIT distance="850" swimtime="00:10:29.08" />
                    <SPLIT distance="900" swimtime="00:11:07.05" />
                    <SPLIT distance="950" swimtime="00:11:44.36" />
                    <SPLIT distance="1000" swimtime="00:12:22.32" />
                    <SPLIT distance="1050" swimtime="00:12:59.43" />
                    <SPLIT distance="1100" swimtime="00:13:37.32" />
                    <SPLIT distance="1150" swimtime="00:14:14.33" />
                    <SPLIT distance="1200" swimtime="00:14:52.24" />
                    <SPLIT distance="1250" swimtime="00:15:29.84" />
                    <SPLIT distance="1300" swimtime="00:16:08.07" />
                    <SPLIT distance="1350" swimtime="00:16:45.49" />
                    <SPLIT distance="1400" swimtime="00:17:23.79" />
                    <SPLIT distance="1450" swimtime="00:18:00.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="458" swimtime="00:00:27.11" resultid="9385" heatid="10623" lane="5" entrytime="00:00:27.51" entrycourse="LCM" />
                <RESULT eventid="1289" points="439" swimtime="00:02:14.17" resultid="9386" heatid="10671" lane="8" entrytime="00:02:15.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.47" />
                    <SPLIT distance="100" swimtime="00:01:05.31" />
                    <SPLIT distance="150" swimtime="00:01:40.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="441" swimtime="00:04:48.91" resultid="9387" heatid="10722" lane="4" entrytime="00:04:41.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                    <SPLIT distance="100" swimtime="00:01:05.60" />
                    <SPLIT distance="150" swimtime="00:01:41.25" />
                    <SPLIT distance="200" swimtime="00:02:18.40" />
                    <SPLIT distance="250" swimtime="00:02:56.04" />
                    <SPLIT distance="300" swimtime="00:03:34.40" />
                    <SPLIT distance="350" swimtime="00:04:12.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kethelyn" lastname="Ribeiro Rodrigues" birthdate="2009-04-24" gender="F" nation="BRA" license="367052" swrid="5600244" athleteid="9124" externalid="367052">
              <RESULTS>
                <RESULT eventid="1095" points="222" swimtime="00:00:40.34" resultid="9125" heatid="10496" lane="7" entrytime="00:00:38.36" entrycourse="LCM" />
                <RESULT eventid="1063" points="255" swimtime="00:03:14.14" resultid="9126" heatid="10470" lane="8" entrytime="00:03:08.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="418" swimtime="00:01:09.13" resultid="9127" heatid="10531" lane="1" entrytime="00:01:07.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="306" swimtime="00:00:39.85" resultid="9128" heatid="10679" lane="0" entrytime="00:00:39.79" entrycourse="LCM" />
                <RESULT eventid="1281" points="426" swimtime="00:02:29.15" resultid="9129" heatid="10657" lane="2" entrytime="00:02:29.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                    <SPLIT distance="100" swimtime="00:01:10.87" />
                    <SPLIT distance="150" swimtime="00:01:49.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="278" swimtime="00:01:27.46" resultid="9130" heatid="10729" lane="0" entrytime="00:01:24.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Inacio Carneiro" birthdate="2009-09-09" gender="M" nation="BRA" license="408023" swrid="5723026" athleteid="9448" externalid="408023">
              <RESULTS>
                <RESULT eventid="1103" points="181" swimtime="00:00:39.31" resultid="9449" heatid="10499" lane="5" />
                <RESULT eventid="1187" points="292" swimtime="00:00:39.09" resultid="9450" heatid="10567" lane="6" />
                <RESULT eventid="1155" points="354" swimtime="00:01:05.59" resultid="9451" heatid="10544" lane="5" entrytime="00:01:05.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="387" swimtime="00:00:28.69" resultid="9452" heatid="10620" lane="4" entrytime="00:00:29.05" entrycourse="LCM" />
                <RESULT eventid="1289" points="331" swimtime="00:02:27.34" resultid="9453" heatid="10667" lane="2" entrytime="00:02:29.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                    <SPLIT distance="100" swimtime="00:01:11.14" />
                    <SPLIT distance="150" swimtime="00:01:50.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="283" swimtime="00:05:35.15" resultid="9454" heatid="10718" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                    <SPLIT distance="100" swimtime="00:01:18.19" />
                    <SPLIT distance="150" swimtime="00:02:00.56" />
                    <SPLIT distance="200" swimtime="00:02:44.38" />
                    <SPLIT distance="250" swimtime="00:03:28.51" />
                    <SPLIT distance="300" swimtime="00:04:13.47" />
                    <SPLIT distance="350" swimtime="00:04:56.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mathias" lastname="Lopes Batista" birthdate="2012-08-22" gender="M" nation="BRA" license="399740" swrid="5652889" athleteid="9258" externalid="399740">
              <RESULTS>
                <RESULT eventid="1071" points="199" swimtime="00:03:11.44" resultid="9259" heatid="10475" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.43" />
                    <SPLIT distance="100" swimtime="00:01:33.82" />
                    <SPLIT distance="150" swimtime="00:02:22.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="248" swimtime="00:01:13.84" resultid="9260" heatid="10540" lane="4" entrytime="00:01:12.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="261" swimtime="00:00:32.69" resultid="9261" heatid="10615" lane="3" entrytime="00:00:32.50" entrycourse="LCM" />
                <RESULT eventid="1305" points="234" swimtime="00:00:38.17" resultid="9262" heatid="10684" lane="8" entrytime="00:00:40.97" entrycourse="LCM" />
                <RESULT eventid="1289" points="207" swimtime="00:02:52.16" resultid="9263" heatid="10665" lane="9" entrytime="00:02:52.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                    <SPLIT distance="100" swimtime="00:01:22.56" />
                    <SPLIT distance="150" swimtime="00:02:07.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="224" swimtime="00:01:24.89" resultid="9264" heatid="10735" lane="5" entrytime="00:01:31.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Nogueira Silva" birthdate="2011-08-13" gender="M" nation="BRA" license="367150" swrid="5588832" athleteid="9166" externalid="367150">
              <RESULTS>
                <RESULT eventid="1087" points="312" swimtime="00:03:04.99" resultid="9167" heatid="10489" lane="6" entrytime="00:03:04.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.77" />
                    <SPLIT distance="100" swimtime="00:01:27.51" />
                    <SPLIT distance="150" swimtime="00:02:16.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="301" swimtime="00:00:38.69" resultid="9168" heatid="10572" lane="7" entrytime="00:00:39.48" entrycourse="LCM" />
                <RESULT eventid="1155" points="398" swimtime="00:01:03.04" resultid="9169" heatid="10545" lane="5" entrytime="00:01:04.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="352" swimtime="00:00:29.61" resultid="9170" heatid="10619" lane="4" entrytime="00:00:29.75" entrycourse="LCM" />
                <RESULT eventid="1219" points="298" swimtime="00:01:25.15" resultid="9171" heatid="10594" lane="4" entrytime="00:01:25.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="329" swimtime="00:02:45.09" resultid="9172" heatid="10647" lane="5" entrytime="00:02:55.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                    <SPLIT distance="100" swimtime="00:01:19.83" />
                    <SPLIT distance="150" swimtime="00:02:08.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Cardim Martins" birthdate="2010-09-01" gender="F" nation="BRA" license="390920" swrid="5600130" athleteid="9305" externalid="390920">
              <RESULTS>
                <RESULT eventid="1095" points="216" swimtime="00:00:40.71" resultid="9306" heatid="10493" lane="5" />
                <RESULT eventid="1063" points="314" swimtime="00:03:01.06" resultid="9307" heatid="10470" lane="4" entrytime="00:02:57.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="359" swimtime="00:01:12.70" resultid="9308" heatid="10527" lane="2" entrytime="00:01:15.44" entrycourse="LCM" />
                <RESULT eventid="1227" points="330" swimtime="00:00:34.14" resultid="9309" heatid="10600" lane="3" />
                <RESULT eventid="1297" points="286" swimtime="00:00:40.74" resultid="9310" heatid="10679" lane="9" entrytime="00:00:39.90" entrycourse="LCM" />
                <RESULT eventid="1365" points="290" swimtime="00:01:26.23" resultid="9311" heatid="10729" lane="1" entrytime="00:01:24.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Gelenski Pelaio" birthdate="2005-10-10" gender="M" nation="BRA" license="281473" swrid="5600173" athleteid="9187" externalid="281473" level="UNIDOMBOSC">
              <RESULTS>
                <RESULT eventid="1155" points="584" swimtime="00:00:55.51" resultid="9188" heatid="10551" lane="1" entrytime="00:00:56.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="563" swimtime="00:00:59.87" resultid="9189" heatid="10711" lane="1" entrytime="00:00:59.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Navarro Silva" birthdate="2011-01-10" gender="F" nation="BRA" license="406711" swrid="5717284" athleteid="9368" externalid="406711">
              <RESULTS>
                <RESULT eventid="1063" points="379" swimtime="00:02:50.12" resultid="9369" heatid="10470" lane="1" entrytime="00:03:06.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="426" swimtime="00:01:08.70" resultid="9370" heatid="10529" lane="5" entrytime="00:01:09.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="422" swimtime="00:00:31.47" resultid="9371" heatid="10605" lane="8" entrytime="00:00:31.50" entrycourse="LCM" />
                <RESULT eventid="1281" points="393" swimtime="00:02:33.09" resultid="9372" heatid="10656" lane="9" entrytime="00:02:36.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                    <SPLIT distance="100" swimtime="00:01:11.97" />
                    <SPLIT distance="150" swimtime="00:01:52.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="332" swimtime="00:05:39.92" resultid="9373" heatid="10713" lane="5" entrytime="00:05:31.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                    <SPLIT distance="100" swimtime="00:01:19.90" />
                    <SPLIT distance="150" swimtime="00:02:03.32" />
                    <SPLIT distance="200" swimtime="00:02:47.25" />
                    <SPLIT distance="250" swimtime="00:03:31.06" />
                    <SPLIT distance="300" swimtime="00:04:15.56" />
                    <SPLIT distance="350" swimtime="00:04:58.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Leticia Durat" birthdate="2008-02-09" gender="F" nation="BRA" license="331636" swrid="5600200" athleteid="9102" externalid="331636">
              <RESULTS>
                <RESULT eventid="1095" points="259" swimtime="00:00:38.31" resultid="9103" heatid="10494" lane="4" />
                <RESULT eventid="1079" points="323" swimtime="00:03:20.42" resultid="9104" heatid="10482" lane="3" entrytime="00:03:21.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.91" />
                    <SPLIT distance="100" swimtime="00:01:35.58" />
                    <SPLIT distance="150" swimtime="00:02:27.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="338" swimtime="00:00:41.83" resultid="9105" heatid="10563" lane="4" entrytime="00:00:40.57" entrycourse="LCM" />
                <RESULT eventid="1147" points="407" swimtime="00:01:09.77" resultid="9106" heatid="10530" lane="7" entrytime="00:01:08.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="333" swimtime="00:01:32.48" resultid="9107" heatid="10585" lane="7" entrytime="00:01:32.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="311" swimtime="00:03:06.09" resultid="9108" heatid="10639" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.89" />
                    <SPLIT distance="100" swimtime="00:01:30.80" />
                    <SPLIT distance="150" swimtime="00:02:22.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juliana" lastname="Moreira Furtado" birthdate="2011-01-27" gender="F" nation="BRA" license="403783" swrid="5684587" athleteid="9279" externalid="403783">
              <RESULTS>
                <RESULT eventid="1095" points="172" swimtime="00:00:43.86" resultid="9280" heatid="10495" lane="2" entrytime="00:00:47.14" entrycourse="LCM" />
                <RESULT eventid="1063" points="217" swimtime="00:03:24.67" resultid="9281" heatid="10469" lane="0">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="312" swimtime="00:01:16.20" resultid="9282" heatid="10527" lane="8" entrytime="00:01:16.91" entrycourse="LCM" />
                <RESULT eventid="1227" points="314" swimtime="00:00:34.72" resultid="9283" heatid="10602" lane="6" entrytime="00:00:35.38" entrycourse="LCM" />
                <RESULT eventid="1281" points="298" swimtime="00:02:48.00" resultid="9284" heatid="10655" lane="0" entrytime="00:02:44.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.36" />
                    <SPLIT distance="100" swimtime="00:01:18.56" />
                    <SPLIT distance="150" swimtime="00:02:03.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="235" swimtime="00:01:32.52" resultid="9285" heatid="10727" lane="1" entrytime="00:01:35.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Prestes Alves Pinto" birthdate="2012-01-19" gender="F" nation="BRA" license="377324" swrid="5588867" athleteid="9238" externalid="377324">
              <RESULTS>
                <RESULT eventid="1095" points="275" swimtime="00:00:37.56" resultid="9239" heatid="10494" lane="8" />
                <RESULT eventid="1063" points="348" swimtime="00:02:54.93" resultid="9240" heatid="10471" lane="1" entrytime="00:02:53.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                    <SPLIT distance="100" swimtime="00:01:23.98" />
                    <SPLIT distance="150" swimtime="00:02:09.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="472" swimtime="00:01:06.37" resultid="9241" heatid="10531" lane="8" entrytime="00:01:07.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="444" swimtime="00:00:30.94" resultid="9242" heatid="10603" lane="4" entrytime="00:00:32.83" entrycourse="LCM" />
                <RESULT eventid="1211" points="277" swimtime="00:01:38.29" resultid="9243" heatid="10583" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="380" swimtime="00:02:54.04" resultid="9244" heatid="10641" lane="9" entrytime="00:03:06.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                    <SPLIT distance="100" swimtime="00:01:20.62" />
                    <SPLIT distance="150" swimtime="00:02:15.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaelle" lastname="Matos De Souza" birthdate="2011-04-24" gender="F" nation="BRA" license="367146" swrid="5628931" athleteid="9152" externalid="367146">
              <RESULTS>
                <RESULT eventid="1063" status="WDR" swimtime="00:00:00.00" resultid="9153" heatid="10470" lane="7" entrytime="00:03:05.29" entrycourse="LCM" />
                <RESULT eventid="1147" status="WDR" swimtime="00:00:00.00" resultid="9154" heatid="10528" lane="3" entrytime="00:01:12.46" entrycourse="LCM" />
                <RESULT eventid="1227" status="WDR" swimtime="00:00:00.00" resultid="9155" heatid="10604" lane="9" entrytime="00:00:32.61" entrycourse="LCM" />
                <RESULT eventid="1297" status="WDR" swimtime="00:00:00.00" resultid="9156" heatid="10676" lane="4" />
                <RESULT eventid="1281" status="WDR" swimtime="00:00:00.00" resultid="9157" heatid="10654" lane="9" />
                <RESULT eventid="1365" status="WDR" swimtime="00:00:00.00" resultid="9158" heatid="10728" lane="6" entrytime="00:01:27.21" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Giulia Aust" birthdate="2011-08-24" gender="F" nation="BRA" license="421352" swrid="4374862" athleteid="9402" externalid="421352">
              <RESULTS>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 19:12)" eventid="1179" status="DSQ" swimtime="00:00:53.97" resultid="9403" heatid="10561" lane="2" />
                <RESULT eventid="1147" points="266" swimtime="00:01:20.35" resultid="9404" heatid="10525" lane="4" entrytime="00:01:20.96" entrycourse="LCM" />
                <RESULT eventid="1227" points="234" swimtime="00:00:38.30" resultid="9405" heatid="10601" lane="3" entrytime="00:00:37.98" entrycourse="LCM" />
                <RESULT eventid="1211" points="156" swimtime="00:01:58.95" resultid="9406" heatid="10583" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="251" swimtime="00:00:42.55" resultid="9407" heatid="10676" lane="3" />
                <RESULT eventid="1365" points="218" swimtime="00:01:34.87" resultid="9408" heatid="10727" lane="8" entrytime="00:01:35.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="16" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1205" points="453" swimtime="00:09:04.80" resultid="9470" heatid="10580" lane="1" entrytime="00:08:46.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.11" />
                    <SPLIT distance="100" swimtime="00:01:01.77" />
                    <SPLIT distance="150" swimtime="00:01:36.05" />
                    <SPLIT distance="200" swimtime="00:02:08.64" />
                    <SPLIT distance="250" swimtime="00:02:38.20" />
                    <SPLIT distance="300" swimtime="00:03:12.66" />
                    <SPLIT distance="350" swimtime="00:03:49.67" />
                    <SPLIT distance="400" swimtime="00:04:26.76" />
                    <SPLIT distance="450" swimtime="00:04:57.29" />
                    <SPLIT distance="500" swimtime="00:05:31.71" />
                    <SPLIT distance="550" swimtime="00:06:09.37" />
                    <SPLIT distance="600" swimtime="00:06:47.50" />
                    <SPLIT distance="650" swimtime="00:07:18.63" />
                    <SPLIT distance="700" swimtime="00:07:54.01" />
                    <SPLIT distance="750" swimtime="00:08:29.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9322" number="1" />
                    <RELAYPOSITION athleteid="9145" number="2" />
                    <RELAYPOSITION athleteid="9291" number="3" />
                    <RELAYPOSITION athleteid="9245" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="19" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1207" points="495" swimtime="00:08:48.97" resultid="9471" heatid="10581" lane="6" entrytime="00:08:16.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.80" />
                    <SPLIT distance="100" swimtime="00:01:01.27" />
                    <SPLIT distance="150" swimtime="00:01:35.44" />
                    <SPLIT distance="200" swimtime="00:02:09.55" />
                    <SPLIT distance="250" swimtime="00:02:37.59" />
                    <SPLIT distance="300" swimtime="00:03:09.82" />
                    <SPLIT distance="350" swimtime="00:03:43.83" />
                    <SPLIT distance="400" swimtime="00:04:17.63" />
                    <SPLIT distance="450" swimtime="00:04:46.01" />
                    <SPLIT distance="500" swimtime="00:05:18.43" />
                    <SPLIT distance="550" swimtime="00:05:54.20" />
                    <SPLIT distance="600" swimtime="00:06:30.05" />
                    <SPLIT distance="650" swimtime="00:07:01.11" />
                    <SPLIT distance="700" swimtime="00:07:34.97" />
                    <SPLIT distance="750" swimtime="00:08:11.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9089" number="1" />
                    <RELAYPOSITION athleteid="9109" number="2" />
                    <RELAYPOSITION athleteid="9395" number="3" />
                    <RELAYPOSITION athleteid="9312" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1203" points="435" swimtime="00:09:12.25" resultid="9472" heatid="10579" lane="3" entrytime="00:09:37.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                    <SPLIT distance="100" swimtime="00:01:05.94" />
                    <SPLIT distance="150" swimtime="00:01:43.47" />
                    <SPLIT distance="200" swimtime="00:02:17.35" />
                    <SPLIT distance="250" swimtime="00:02:47.47" />
                    <SPLIT distance="300" swimtime="00:03:23.02" />
                    <SPLIT distance="350" swimtime="00:03:58.92" />
                    <SPLIT distance="400" swimtime="00:04:33.35" />
                    <SPLIT distance="450" swimtime="00:05:05.43" />
                    <SPLIT distance="500" swimtime="00:05:40.43" />
                    <SPLIT distance="550" swimtime="00:06:15.71" />
                    <SPLIT distance="600" swimtime="00:06:51.56" />
                    <SPLIT distance="650" swimtime="00:07:22.15" />
                    <SPLIT distance="700" swimtime="00:07:56.82" />
                    <SPLIT distance="750" swimtime="00:08:34.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9272" number="1" />
                    <RELAYPOSITION athleteid="9138" number="2" />
                    <RELAYPOSITION athleteid="9197" number="3" />
                    <RELAYPOSITION athleteid="9204" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1331" points="505" swimtime="00:04:19.55" resultid="9473" heatid="10698" lane="3" entrytime="00:04:14.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                    <SPLIT distance="150" swimtime="00:01:40.56" />
                    <SPLIT distance="200" swimtime="00:02:21.79" />
                    <SPLIT distance="250" swimtime="00:02:50.74" />
                    <SPLIT distance="300" swimtime="00:03:24.22" />
                    <SPLIT distance="350" swimtime="00:03:50.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9115" number="1" />
                    <RELAYPOSITION athleteid="9381" number="2" />
                    <RELAYPOSITION athleteid="9118" number="3" />
                    <RELAYPOSITION athleteid="9109" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1399" points="600" swimtime="00:03:43.07" resultid="9478" heatid="10753" lane="5" entrytime="00:03:41.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.49" />
                    <SPLIT distance="100" swimtime="00:00:55.86" />
                    <SPLIT distance="150" swimtime="00:01:21.63" />
                    <SPLIT distance="200" swimtime="00:01:49.71" />
                    <SPLIT distance="250" swimtime="00:02:16.96" />
                    <SPLIT distance="300" swimtime="00:02:47.55" />
                    <SPLIT distance="350" swimtime="00:03:13.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9187" number="1" />
                    <RELAYPOSITION athleteid="9118" number="2" />
                    <RELAYPOSITION athleteid="9089" number="3" />
                    <RELAYPOSITION athleteid="9109" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1329" points="314" swimtime="00:05:04.19" resultid="9474" heatid="10697" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                    <SPLIT distance="100" swimtime="00:01:16.09" />
                    <SPLIT distance="150" swimtime="00:01:55.61" />
                    <SPLIT distance="200" swimtime="00:02:43.85" />
                    <SPLIT distance="250" swimtime="00:03:17.95" />
                    <SPLIT distance="300" swimtime="00:04:00.98" />
                    <SPLIT distance="350" swimtime="00:04:30.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9291" number="1" />
                    <RELAYPOSITION athleteid="9448" number="2" />
                    <RELAYPOSITION athleteid="9455" number="3" />
                    <RELAYPOSITION athleteid="9438" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1397" status="DNS" swimtime="00:00:00.00" resultid="9479" heatid="10752" lane="2">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9291" number="1" />
                    <RELAYPOSITION athleteid="9448" number="2" />
                    <RELAYPOSITION athleteid="9438" number="3" />
                    <RELAYPOSITION athleteid="9388" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1323" points="231" swimtime="00:05:36.90" resultid="9475" heatid="10693" lane="5" entrytime="00:04:51.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                    <SPLIT distance="100" swimtime="00:01:26.67" />
                    <SPLIT distance="150" swimtime="00:02:06.47" />
                    <SPLIT distance="200" swimtime="00:02:54.11" />
                    <SPLIT distance="250" swimtime="00:03:30.60" />
                    <SPLIT distance="300" swimtime="00:04:18.76" />
                    <SPLIT distance="350" swimtime="00:04:54.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9258" number="1" />
                    <RELAYPOSITION athleteid="9190" number="2" />
                    <RELAYPOSITION athleteid="9341" number="3" />
                    <RELAYPOSITION athleteid="9252" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1391" status="WDR" swimtime="00:00:00.00" resultid="9482" heatid="10748" lane="4" entrytime="00:04:15.70">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9252" number="1" />
                    <RELAYPOSITION athleteid="9258" number="2" />
                    <RELAYPOSITION athleteid="9341" number="3" />
                    <RELAYPOSITION athleteid="9190" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 19:52)" eventid="1327" status="DSQ" swimtime="00:05:15.14" resultid="9476" heatid="10696" lane="5" entrytime="00:04:25.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.75" />
                    <SPLIT distance="150" swimtime="00:02:08.06" />
                    <SPLIT distance="200" swimtime="00:02:55.37" />
                    <SPLIT distance="250" swimtime="00:03:29.21" />
                    <SPLIT distance="300" swimtime="00:04:04.94" />
                    <SPLIT distance="350" swimtime="00:04:38.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9415" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="9388" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="9245" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="9442" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1395" points="476" swimtime="00:04:01.02" resultid="9480" heatid="10751" lane="3" entrytime="00:03:56.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                    <SPLIT distance="100" swimtime="00:00:58.29" />
                    <SPLIT distance="150" swimtime="00:01:27.50" />
                    <SPLIT distance="200" swimtime="00:02:00.72" />
                    <SPLIT distance="250" swimtime="00:02:29.06" />
                    <SPLIT distance="300" swimtime="00:03:00.56" />
                    <SPLIT distance="350" swimtime="00:03:29.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9322" number="1" />
                    <RELAYPOSITION athleteid="9173" number="2" />
                    <RELAYPOSITION athleteid="9145" number="3" />
                    <RELAYPOSITION athleteid="9245" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1325" points="437" swimtime="00:04:32.45" resultid="9477" heatid="10695" lane="3" entrytime="00:04:50.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                    <SPLIT distance="100" swimtime="00:01:08.79" />
                    <SPLIT distance="150" swimtime="00:01:44.14" />
                    <SPLIT distance="200" swimtime="00:02:27.15" />
                    <SPLIT distance="250" swimtime="00:02:56.04" />
                    <SPLIT distance="300" swimtime="00:03:30.33" />
                    <SPLIT distance="350" swimtime="00:03:59.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9138" number="1" />
                    <RELAYPOSITION athleteid="9159" number="2" />
                    <RELAYPOSITION athleteid="9272" number="3" />
                    <RELAYPOSITION athleteid="9166" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1393" points="427" swimtime="00:04:09.80" resultid="9481" heatid="10750" lane="6" entrytime="00:04:15.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.54" />
                    <SPLIT distance="100" swimtime="00:01:00.98" />
                    <SPLIT distance="150" swimtime="00:01:30.97" />
                    <SPLIT distance="200" swimtime="00:02:04.07" />
                    <SPLIT distance="250" swimtime="00:02:33.84" />
                    <SPLIT distance="300" swimtime="00:03:06.54" />
                    <SPLIT distance="350" swimtime="00:03:36.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9272" number="1" />
                    <RELAYPOSITION athleteid="9138" number="2" />
                    <RELAYPOSITION athleteid="9166" number="3" />
                    <RELAYPOSITION athleteid="9204" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1327" points="427" swimtime="00:04:34.56" resultid="9488" heatid="10696" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                    <SPLIT distance="100" swimtime="00:01:17.75" />
                    <SPLIT distance="150" swimtime="00:01:51.63" />
                    <SPLIT distance="200" swimtime="00:02:30.79" />
                    <SPLIT distance="250" swimtime="00:03:00.52" />
                    <SPLIT distance="300" swimtime="00:03:36.89" />
                    <SPLIT distance="350" swimtime="00:04:04.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9334" number="1" />
                    <RELAYPOSITION athleteid="9173" number="2" />
                    <RELAYPOSITION athleteid="9145" number="3" />
                    <RELAYPOSITION athleteid="9322" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1395" points="340" swimtime="00:04:29.51" resultid="9490" heatid="10751" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="150" swimtime="00:01:37.94" />
                    <SPLIT distance="200" swimtime="00:02:13.68" />
                    <SPLIT distance="250" swimtime="00:02:48.65" />
                    <SPLIT distance="300" swimtime="00:03:24.75" />
                    <SPLIT distance="350" swimtime="00:03:55.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9455" number="1" />
                    <RELAYPOSITION athleteid="9415" number="2" />
                    <RELAYPOSITION athleteid="9442" number="3" />
                    <RELAYPOSITION athleteid="9334" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1325" points="275" swimtime="00:05:17.65" resultid="9489" heatid="10694" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.47" />
                    <SPLIT distance="100" swimtime="00:01:23.82" />
                    <SPLIT distance="150" swimtime="00:02:08.44" />
                    <SPLIT distance="200" swimtime="00:02:56.50" />
                    <SPLIT distance="250" swimtime="00:03:29.32" />
                    <SPLIT distance="300" swimtime="00:04:07.04" />
                    <SPLIT distance="350" swimtime="00:04:40.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9204" number="1" />
                    <RELAYPOSITION athleteid="9348" number="2" />
                    <RELAYPOSITION athleteid="9197" number="3" />
                    <RELAYPOSITION athleteid="9374" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1393" points="321" swimtime="00:04:34.88" resultid="9491" heatid="10750" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                    <SPLIT distance="100" swimtime="00:01:11.58" />
                    <SPLIT distance="150" swimtime="00:01:46.73" />
                    <SPLIT distance="200" swimtime="00:02:25.73" />
                    <SPLIT distance="250" swimtime="00:02:56.44" />
                    <SPLIT distance="300" swimtime="00:03:31.99" />
                    <SPLIT distance="350" swimtime="00:04:02.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9374" number="1" />
                    <RELAYPOSITION athleteid="9348" number="2" />
                    <RELAYPOSITION athleteid="9159" number="3" />
                    <RELAYPOSITION athleteid="9197" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="F" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1197" points="412" swimtime="00:10:14.42" resultid="9462" heatid="10577" lane="7" entrytime="00:09:37.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                    <SPLIT distance="100" swimtime="00:01:11.66" />
                    <SPLIT distance="150" swimtime="00:01:50.98" />
                    <SPLIT distance="200" swimtime="00:02:28.66" />
                    <SPLIT distance="250" swimtime="00:03:01.82" />
                    <SPLIT distance="300" swimtime="00:03:41.60" />
                    <SPLIT distance="350" swimtime="00:04:23.66" />
                    <SPLIT distance="400" swimtime="00:05:03.30" />
                    <SPLIT distance="450" swimtime="00:05:37.47" />
                    <SPLIT distance="500" swimtime="00:06:17.40" />
                    <SPLIT distance="550" swimtime="00:06:59.56" />
                    <SPLIT distance="600" swimtime="00:07:39.58" />
                    <SPLIT distance="650" swimtime="00:08:14.47" />
                    <SPLIT distance="700" swimtime="00:08:53.12" />
                    <SPLIT distance="750" swimtime="00:09:33.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9217" number="1" />
                    <RELAYPOSITION athleteid="9180" number="2" />
                    <RELAYPOSITION athleteid="9231" number="3" />
                    <RELAYPOSITION athleteid="9298" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1195" points="407" swimtime="00:10:16.98" resultid="9463" heatid="10576" lane="1" entrytime="00:10:00.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                    <SPLIT distance="100" swimtime="00:01:12.57" />
                    <SPLIT distance="150" swimtime="00:01:51.98" />
                    <SPLIT distance="200" swimtime="00:02:29.24" />
                    <SPLIT distance="250" swimtime="00:03:03.98" />
                    <SPLIT distance="300" swimtime="00:03:43.66" />
                    <SPLIT distance="350" swimtime="00:04:22.93" />
                    <SPLIT distance="400" swimtime="00:05:00.57" />
                    <SPLIT distance="450" swimtime="00:05:35.69" />
                    <SPLIT distance="500" swimtime="00:06:14.29" />
                    <SPLIT distance="550" swimtime="00:06:55.03" />
                    <SPLIT distance="600" swimtime="00:07:35.30" />
                    <SPLIT distance="650" swimtime="00:08:10.92" />
                    <SPLIT distance="700" swimtime="00:08:52.91" />
                    <SPLIT distance="750" swimtime="00:09:35.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9238" number="1" />
                    <RELAYPOSITION athleteid="9265" number="2" />
                    <RELAYPOSITION athleteid="9368" number="3" />
                    <RELAYPOSITION athleteid="9426" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1315" points="231" swimtime="00:06:13.85" resultid="9464" heatid="10689" lane="4" entrytime="00:05:17.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.97" />
                    <SPLIT distance="100" swimtime="00:01:31.49" />
                    <SPLIT distance="150" swimtime="00:02:14.84" />
                    <SPLIT distance="200" swimtime="00:03:03.71" />
                    <SPLIT distance="250" swimtime="00:03:49.00" />
                    <SPLIT distance="350" swimtime="00:05:28.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9279" number="1" />
                    <RELAYPOSITION athleteid="9131" number="2" />
                    <RELAYPOSITION athleteid="9368" number="3" />
                    <RELAYPOSITION athleteid="9402" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1383" points="335" swimtime="00:04:59.25" resultid="9469" heatid="10744" lane="6" entrytime="00:04:34.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                    <SPLIT distance="100" swimtime="00:01:22.56" />
                    <SPLIT distance="150" swimtime="00:01:58.06" />
                    <SPLIT distance="200" swimtime="00:02:38.51" />
                    <SPLIT distance="250" swimtime="00:03:12.69" />
                    <SPLIT distance="300" swimtime="00:03:51.31" />
                    <SPLIT distance="350" swimtime="00:04:24.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9402" number="1" />
                    <RELAYPOSITION athleteid="9279" number="2" />
                    <RELAYPOSITION athleteid="9131" number="3" />
                    <RELAYPOSITION athleteid="9368" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="F" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1317" points="400" swimtime="00:05:11.40" resultid="9465" heatid="10690" lane="2" entrytime="00:05:10.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.74" />
                    <SPLIT distance="100" swimtime="00:01:25.98" />
                    <SPLIT distance="150" swimtime="00:02:05.27" />
                    <SPLIT distance="200" swimtime="00:02:48.56" />
                    <SPLIT distance="250" swimtime="00:03:23.74" />
                    <SPLIT distance="300" swimtime="00:04:04.19" />
                    <SPLIT distance="350" swimtime="00:04:35.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9305" number="1" />
                    <RELAYPOSITION athleteid="9217" number="2" />
                    <RELAYPOSITION athleteid="9180" number="3" />
                    <RELAYPOSITION athleteid="9298" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1385" points="438" swimtime="00:04:33.79" resultid="9468" heatid="10745" lane="2" entrytime="00:04:16.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.66" />
                    <SPLIT distance="100" swimtime="00:01:07.77" />
                    <SPLIT distance="150" swimtime="00:01:40.15" />
                    <SPLIT distance="200" swimtime="00:02:16.35" />
                    <SPLIT distance="250" swimtime="00:02:49.51" />
                    <SPLIT distance="300" swimtime="00:03:26.82" />
                    <SPLIT distance="350" swimtime="00:03:58.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9180" number="1" />
                    <RELAYPOSITION athleteid="9217" number="2" />
                    <RELAYPOSITION athleteid="9231" number="3" />
                    <RELAYPOSITION athleteid="9298" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1313" points="363" swimtime="00:05:21.89" resultid="9466" heatid="10688" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.42" />
                    <SPLIT distance="100" swimtime="00:01:19.45" />
                    <SPLIT distance="150" swimtime="00:02:02.97" />
                    <SPLIT distance="200" swimtime="00:02:55.29" />
                    <SPLIT distance="250" swimtime="00:03:31.54" />
                    <SPLIT distance="300" swimtime="00:04:15.83" />
                    <SPLIT distance="350" swimtime="00:04:46.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9426" number="1" />
                    <RELAYPOSITION athleteid="9210" number="2" />
                    <RELAYPOSITION athleteid="9265" number="3" />
                    <RELAYPOSITION athleteid="9238" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" points="412" swimtime="00:04:39.39" resultid="9467" heatid="10743" lane="3" entrytime="00:05:30.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                    <SPLIT distance="100" swimtime="00:01:15.93" />
                    <SPLIT distance="150" swimtime="00:01:50.76" />
                    <SPLIT distance="200" swimtime="00:02:27.91" />
                    <SPLIT distance="250" swimtime="00:02:58.83" />
                    <SPLIT distance="300" swimtime="00:03:33.66" />
                    <SPLIT distance="350" swimtime="00:04:05.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9210" number="1" />
                    <RELAYPOSITION athleteid="9426" number="2" />
                    <RELAYPOSITION athleteid="9238" number="3" />
                    <RELAYPOSITION athleteid="9265" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1113" points="407" swimtime="00:04:53.34" resultid="9483" heatid="10510" lane="2" entrytime="00:04:53.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                    <SPLIT distance="100" swimtime="00:01:09.44" />
                    <SPLIT distance="150" swimtime="00:01:53.03" />
                    <SPLIT distance="200" swimtime="00:02:40.81" />
                    <SPLIT distance="250" swimtime="00:03:09.94" />
                    <SPLIT distance="300" swimtime="00:03:44.85" />
                    <SPLIT distance="350" swimtime="00:04:18.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9138" number="1" />
                    <RELAYPOSITION athleteid="9131" number="2" />
                    <RELAYPOSITION athleteid="9272" number="3" />
                    <RELAYPOSITION athleteid="9368" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1111" points="321" swimtime="00:05:17.50" resultid="9484" heatid="10509" lane="6" entrytime="00:05:06.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.67" />
                    <SPLIT distance="100" swimtime="00:01:21.77" />
                    <SPLIT distance="150" swimtime="00:02:00.67" />
                    <SPLIT distance="200" swimtime="00:02:47.04" />
                    <SPLIT distance="250" swimtime="00:03:21.60" />
                    <SPLIT distance="300" swimtime="00:04:05.17" />
                    <SPLIT distance="350" swimtime="00:04:37.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9238" number="1" />
                    <RELAYPOSITION athleteid="9190" number="2" />
                    <RELAYPOSITION athleteid="9265" number="3" />
                    <RELAYPOSITION athleteid="9258" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1247" points="443" swimtime="00:04:45.18" resultid="9485" heatid="10631" lane="3" entrytime="00:04:33.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                    <SPLIT distance="100" swimtime="00:01:04.57" />
                    <SPLIT distance="150" swimtime="00:01:46.78" />
                    <SPLIT distance="200" swimtime="00:02:37.10" />
                    <SPLIT distance="250" swimtime="00:03:07.61" />
                    <SPLIT distance="300" swimtime="00:03:42.22" />
                    <SPLIT distance="350" swimtime="00:04:12.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9118" number="1" />
                    <RELAYPOSITION athleteid="9102" number="2" />
                    <RELAYPOSITION athleteid="9089" number="3" />
                    <RELAYPOSITION athleteid="9082" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1243" points="420" swimtime="00:04:50.11" resultid="9486" heatid="10629" lane="5" entrytime="00:04:31.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                    <SPLIT distance="100" swimtime="00:01:16.28" />
                    <SPLIT distance="150" swimtime="00:01:55.80" />
                    <SPLIT distance="200" swimtime="00:02:38.94" />
                    <SPLIT distance="250" swimtime="00:03:08.08" />
                    <SPLIT distance="300" swimtime="00:03:44.46" />
                    <SPLIT distance="350" swimtime="00:04:15.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9334" number="1" />
                    <RELAYPOSITION athleteid="9217" number="2" />
                    <RELAYPOSITION athleteid="9145" number="3" />
                    <RELAYPOSITION athleteid="9180" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1245" points="341" swimtime="00:05:11.03" resultid="9487" heatid="10630" lane="2" entrytime="00:05:03.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.41" />
                    <SPLIT distance="100" swimtime="00:01:26.53" />
                    <SPLIT distance="150" swimtime="00:02:07.53" />
                    <SPLIT distance="200" swimtime="00:02:56.09" />
                    <SPLIT distance="250" swimtime="00:03:30.85" />
                    <SPLIT distance="300" swimtime="00:04:07.78" />
                    <SPLIT distance="350" swimtime="00:04:37.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9124" number="1" />
                    <RELAYPOSITION athleteid="9231" number="2" />
                    <RELAYPOSITION athleteid="9245" number="3" />
                    <RELAYPOSITION athleteid="9438" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 12:08), Na volta dos 250m (Borboleta, Revezamento Medley)." eventid="1113" status="DSQ" swimtime="00:05:27.61" resultid="9492" heatid="10510" lane="7" entrytime="00:05:15.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.89" />
                    <SPLIT distance="100" swimtime="00:01:33.65" />
                    <SPLIT distance="150" swimtime="00:02:10.65" />
                    <SPLIT distance="200" swimtime="00:02:54.39" />
                    <SPLIT distance="250" swimtime="00:03:26.29" />
                    <SPLIT distance="300" swimtime="00:04:03.96" />
                    <SPLIT distance="350" swimtime="00:04:44.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9279" number="1" />
                    <RELAYPOSITION athleteid="9159" number="2" />
                    <RELAYPOSITION athleteid="9197" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="9286" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1111" points="274" swimtime="00:05:34.53" resultid="9493" heatid="10509" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                    <SPLIT distance="100" swimtime="00:01:20.28" />
                    <SPLIT distance="150" swimtime="00:02:03.88" />
                    <SPLIT distance="200" swimtime="00:02:53.34" />
                    <SPLIT distance="250" swimtime="00:03:28.35" />
                    <SPLIT distance="300" swimtime="00:04:16.37" />
                    <SPLIT distance="350" swimtime="00:04:51.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9426" number="1" />
                    <RELAYPOSITION athleteid="9210" number="2" />
                    <RELAYPOSITION athleteid="9341" number="3" />
                    <RELAYPOSITION athleteid="9252" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1243" points="367" swimtime="00:05:03.49" resultid="9494" heatid="10629" lane="3" entrytime="00:04:35.37">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9305" number="1" />
                    <RELAYPOSITION athleteid="9173" number="2" />
                    <RELAYPOSITION athleteid="9298" number="3" />
                    <RELAYPOSITION athleteid="9322" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="439" nation="BRA" region="RJ" clubid="8830" swrid="75483" name="Fluminense Football Club" shortname="Ffc/Rj">
          <ATHLETES>
            <ATHLETE firstname="Felipe" lastname="Chi Kravchychyn" birthdate="2009-09-27" gender="M" nation="BRA" license="344268" swrid="5600134" athleteid="8831" externalid="344268">
              <RESULTS>
                <RESULT eventid="1087" points="622" status="EXH" swimtime="00:02:26.96" resultid="8832" heatid="10492" lane="5" entrytime="00:02:26.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                    <SPLIT distance="100" swimtime="00:01:10.77" />
                    <SPLIT distance="150" swimtime="00:01:49.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="451" status="EXH" swimtime="00:02:25.91" resultid="8833" heatid="10479" lane="9" entrytime="00:02:27.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                    <SPLIT distance="100" swimtime="00:01:10.06" />
                    <SPLIT distance="150" swimtime="00:01:48.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="438" status="EXH" swimtime="00:02:25.22" resultid="8834" heatid="10558" lane="8" entrytime="00:02:23.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                    <SPLIT distance="100" swimtime="00:01:06.11" />
                    <SPLIT distance="150" swimtime="00:01:44.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="573" status="EXH" swimtime="00:04:51.82" resultid="8835" heatid="10523" lane="5" entrytime="00:04:49.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                    <SPLIT distance="100" swimtime="00:01:05.42" />
                    <SPLIT distance="150" swimtime="00:01:44.75" />
                    <SPLIT distance="200" swimtime="00:02:23.48" />
                    <SPLIT distance="250" swimtime="00:03:03.58" />
                    <SPLIT distance="300" swimtime="00:03:43.47" />
                    <SPLIT distance="350" swimtime="00:04:18.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="533" status="EXH" swimtime="00:17:53.59" resultid="8836" heatid="10638" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                    <SPLIT distance="100" swimtime="00:01:05.21" />
                    <SPLIT distance="150" swimtime="00:01:40.77" />
                    <SPLIT distance="200" swimtime="00:02:16.98" />
                    <SPLIT distance="250" swimtime="00:02:52.72" />
                    <SPLIT distance="300" swimtime="00:03:28.95" />
                    <SPLIT distance="350" swimtime="00:04:04.23" />
                    <SPLIT distance="400" swimtime="00:04:40.53" />
                    <SPLIT distance="450" swimtime="00:05:16.51" />
                    <SPLIT distance="500" swimtime="00:05:53.01" />
                    <SPLIT distance="550" swimtime="00:06:28.89" />
                    <SPLIT distance="600" swimtime="00:07:05.17" />
                    <SPLIT distance="650" swimtime="00:07:40.81" />
                    <SPLIT distance="700" swimtime="00:08:16.94" />
                    <SPLIT distance="750" swimtime="00:08:52.75" />
                    <SPLIT distance="800" swimtime="00:09:28.67" />
                    <SPLIT distance="850" swimtime="00:10:04.73" />
                    <SPLIT distance="900" swimtime="00:10:41.01" />
                    <SPLIT distance="950" swimtime="00:11:16.90" />
                    <SPLIT distance="1000" swimtime="00:11:53.09" />
                    <SPLIT distance="1050" swimtime="00:12:29.05" />
                    <SPLIT distance="1100" swimtime="00:13:05.43" />
                    <SPLIT distance="1150" swimtime="00:13:41.72" />
                    <SPLIT distance="1200" swimtime="00:14:18.21" />
                    <SPLIT distance="1250" swimtime="00:14:54.48" />
                    <SPLIT distance="1300" swimtime="00:15:30.91" />
                    <SPLIT distance="1350" swimtime="00:16:07.43" />
                    <SPLIT distance="1400" swimtime="00:16:44.12" />
                    <SPLIT distance="1450" swimtime="00:17:19.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="545" status="EXH" swimtime="00:02:04.80" resultid="8837" heatid="10661" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.14" />
                    <SPLIT distance="100" swimtime="00:00:59.59" />
                    <SPLIT distance="150" swimtime="00:01:32.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3501" nation="BRA" region="PR" clubid="7189" swrid="93752" name="Ortega &amp; De Souza Jesus" shortname="Aquafoz">
          <ATHLETES>
            <ATHLETE firstname="Julia" lastname="Victoria Portela" birthdate="2009-12-04" gender="F" nation="BRA" license="383047" swrid="5596945" athleteid="7214" externalid="383047">
              <RESULTS>
                <RESULT eventid="1147" points="480" swimtime="00:01:06.02" resultid="7215" heatid="10533" lane="0" entrytime="00:01:05.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="496" swimtime="00:00:29.82" resultid="7216" heatid="10609" lane="1" entrytime="00:00:29.11" entrycourse="LCM" />
                <RESULT eventid="1281" points="397" swimtime="00:02:32.58" resultid="7217" heatid="10656" lane="4" entrytime="00:02:30.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                    <SPLIT distance="100" swimtime="00:01:10.56" />
                    <SPLIT distance="150" swimtime="00:01:51.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulo" lastname="Antonio Sousa" birthdate="2012-03-17" gender="M" nation="BRA" license="407497" swrid="5721498" athleteid="7250" externalid="407497">
              <RESULTS>
                <RESULT eventid="1103" points="135" swimtime="00:00:43.35" resultid="7251" heatid="10500" lane="8" />
                <RESULT eventid="1187" points="234" swimtime="00:00:42.07" resultid="7252" heatid="10569" lane="4" />
                <RESULT eventid="1155" points="253" swimtime="00:01:13.28" resultid="7253" heatid="10535" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="239" swimtime="00:00:33.69" resultid="7254" heatid="10610" lane="4" />
                <RESULT eventid="1305" points="173" swimtime="00:00:42.25" resultid="7255" heatid="10682" lane="0" />
                <RESULT eventid="1373" points="201" swimtime="00:01:28.00" resultid="7256" heatid="10735" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Gustavo Cunha" birthdate="2011-01-31" gender="M" nation="BRA" license="392836" swrid="5641764" athleteid="7238" externalid="392836">
              <RESULTS>
                <RESULT eventid="1155" points="296" swimtime="00:01:09.61" resultid="7239" heatid="10541" lane="7" entrytime="00:01:11.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="326" swimtime="00:00:30.36" resultid="7240" heatid="10615" lane="8" entrytime="00:00:33.08" entrycourse="LCM" />
                <RESULT eventid="1305" points="239" swimtime="00:00:37.93" resultid="7241" heatid="10681" lane="6" />
                <RESULT eventid="1373" points="205" swimtime="00:01:27.38" resultid="7242" heatid="10733" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julio" lastname="Heck" birthdate="1998-02-15" gender="M" nation="BRA" license="185880" swrid="5596906" athleteid="7204" externalid="185880">
              <RESULTS>
                <RESULT eventid="1103" points="509" swimtime="00:00:27.89" resultid="7205" heatid="10508" lane="1" entrytime="00:00:27.44" entrycourse="LCM" />
                <RESULT eventid="1155" points="634" swimtime="00:00:54.00" resultid="7206" heatid="10552" lane="2" entrytime="00:00:53.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="636" swimtime="00:00:24.31" resultid="7207" heatid="10628" lane="7" entrytime="00:00:24.41" entrycourse="LCM" />
                <RESULT eventid="1305" points="444" swimtime="00:00:30.86" resultid="7208" heatid="10686" lane="7" entrytime="00:00:31.55" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luisa" lastname="Franco" birthdate="2010-06-09" gender="F" nation="BRA" license="383849" swrid="5596896" athleteid="7194" externalid="383849">
              <RESULTS>
                <RESULT eventid="1095" points="431" swimtime="00:00:32.33" resultid="7195" heatid="10496" lane="5" entrytime="00:00:36.53" entrycourse="LCM" />
                <RESULT eventid="1227" points="438" swimtime="00:00:31.08" resultid="7196" heatid="10604" lane="1" entrytime="00:00:32.23" entrycourse="LCM" />
                <RESULT eventid="1281" points="428" swimtime="00:02:28.82" resultid="7197" heatid="10656" lane="7" entrytime="00:02:33.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                    <SPLIT distance="100" swimtime="00:01:11.81" />
                    <SPLIT distance="150" swimtime="00:01:51.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="406" swimtime="00:01:14.49" resultid="7198" heatid="10699" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Geórgia" lastname="Adeli Jesus" birthdate="2008-03-27" gender="F" nation="BRA" license="312649" swrid="5596864" athleteid="7209" externalid="312649">
              <RESULTS>
                <RESULT eventid="1147" points="432" swimtime="00:01:08.40" resultid="7210" heatid="10529" lane="3" entrytime="00:01:10.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="370" swimtime="00:11:14.76" resultid="7211" heatid="10633" lane="3" entrytime="00:11:10.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.17" />
                    <SPLIT distance="100" swimtime="00:01:11.71" />
                    <SPLIT distance="150" swimtime="00:01:50.78" />
                    <SPLIT distance="200" swimtime="00:02:33.05" />
                    <SPLIT distance="250" swimtime="00:03:14.96" />
                    <SPLIT distance="300" swimtime="00:03:58.47" />
                    <SPLIT distance="350" swimtime="00:04:41.88" />
                    <SPLIT distance="400" swimtime="00:05:26.67" />
                    <SPLIT distance="450" swimtime="00:06:11.01" />
                    <SPLIT distance="500" swimtime="00:06:57.57" />
                    <SPLIT distance="550" swimtime="00:07:41.38" />
                    <SPLIT distance="600" swimtime="00:08:25.66" />
                    <SPLIT distance="650" swimtime="00:09:09.49" />
                    <SPLIT distance="700" swimtime="00:09:52.05" />
                    <SPLIT distance="750" swimtime="00:10:33.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="426" swimtime="00:02:29.14" resultid="7212" heatid="10657" lane="5" entrytime="00:02:28.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                    <SPLIT distance="100" swimtime="00:01:09.88" />
                    <SPLIT distance="150" swimtime="00:01:49.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="347" swimtime="00:05:34.74" resultid="7213" heatid="10714" lane="2" entrytime="00:05:18.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="100" swimtime="00:01:13.94" />
                    <SPLIT distance="150" swimtime="00:01:55.70" />
                    <SPLIT distance="200" swimtime="00:02:39.01" />
                    <SPLIT distance="250" swimtime="00:03:22.36" />
                    <SPLIT distance="300" swimtime="00:04:06.97" />
                    <SPLIT distance="350" swimtime="00:04:51.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Afonso Proteti" birthdate="2002-03-19" gender="M" nation="BRA" license="190464" swrid="5596865" athleteid="7199" externalid="190464">
              <RESULTS>
                <RESULT eventid="1103" points="624" swimtime="00:00:26.06" resultid="7200" heatid="10508" lane="5" entrytime="00:00:25.19" entrycourse="LCM" />
                <RESULT eventid="1187" points="537" swimtime="00:00:31.91" resultid="7201" heatid="10566" lane="5" />
                <RESULT eventid="1305" points="561" swimtime="00:00:28.54" resultid="7202" heatid="10687" lane="5" entrytime="00:00:28.62" entrycourse="LCM" />
                <RESULT eventid="1341" points="613" swimtime="00:00:58.20" resultid="7203" heatid="10711" lane="5" entrytime="00:00:57.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="Wirtti" birthdate="2011-01-14" gender="M" nation="BRA" license="383854" swrid="4917570" athleteid="7228" externalid="383854">
              <RESULTS>
                <RESULT eventid="1103" points="320" swimtime="00:00:32.53" resultid="7229" heatid="10503" lane="4" entrytime="00:00:34.80" entrycourse="LCM" />
                <RESULT eventid="1155" points="384" swimtime="00:01:03.80" resultid="7230" heatid="10545" lane="9" entrytime="00:01:05.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="395" swimtime="00:00:28.48" resultid="7231" heatid="10620" lane="0" entrytime="00:00:29.65" entrycourse="LCM" />
                <RESULT eventid="1305" points="332" swimtime="00:00:33.98" resultid="7232" heatid="10685" lane="0" entrytime="00:00:35.53" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Marques Lima" birthdate="2010-04-30" gender="F" nation="BRA" license="383051" swrid="5596913" athleteid="7218" externalid="383051">
              <RESULTS>
                <RESULT eventid="1063" points="350" swimtime="00:02:54.63" resultid="7219" heatid="10470" lane="3" entrytime="00:02:57.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="371" swimtime="00:00:32.85" resultid="7220" heatid="10603" lane="5" entrytime="00:00:32.86" entrycourse="LCM" />
                <RESULT eventid="1297" points="404" swimtime="00:00:36.32" resultid="7221" heatid="10679" lane="6" entrytime="00:00:37.89" entrycourse="LCM" />
                <RESULT eventid="1365" points="371" swimtime="00:01:19.46" resultid="7222" heatid="10729" lane="3" entrytime="00:01:22.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kauan" lastname="Matheus Cunha" birthdate="2011-01-31" gender="M" nation="BRA" license="392834" swrid="5641770" athleteid="7233" externalid="392834">
              <RESULTS>
                <RESULT eventid="1103" points="217" swimtime="00:00:37.04" resultid="7234" heatid="10503" lane="8" entrytime="00:00:36.88" entrycourse="LCM" />
                <RESULT eventid="1155" points="256" swimtime="00:01:13.06" resultid="7235" heatid="10540" lane="0" entrytime="00:01:13.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="273" swimtime="00:00:32.21" resultid="7236" heatid="10616" lane="0" entrytime="00:00:32.21" entrycourse="LCM" />
                <RESULT eventid="1341" points="184" swimtime="00:01:26.84" resultid="7237" heatid="10705" lane="0" entrytime="00:01:38.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Gabriel Serighelli" birthdate="1999-03-12" gender="M" nation="BRA" license="121253" swrid="5596899" athleteid="7190" externalid="121253">
              <RESULTS>
                <RESULT eventid="1235" points="526" swimtime="00:00:25.89" resultid="7191" heatid="10627" lane="0" entrytime="00:00:25.40" entrycourse="LCM" />
                <RESULT eventid="1305" points="524" swimtime="00:00:29.21" resultid="7192" heatid="10687" lane="3" entrytime="00:00:29.08" entrycourse="LCM" />
                <RESULT eventid="1373" points="459" swimtime="00:01:06.86" resultid="7193" heatid="10741" lane="8" entrytime="00:01:06.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Xavier" birthdate="2011-10-14" gender="M" nation="BRA" license="370564" swrid="5596949" athleteid="7223" externalid="370564">
              <RESULTS>
                <RESULT eventid="1087" points="300" swimtime="00:03:07.25" resultid="7224" heatid="10489" lane="9" entrytime="00:03:12.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.26" />
                    <SPLIT distance="100" swimtime="00:01:29.31" />
                    <SPLIT distance="150" swimtime="00:02:17.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="263" swimtime="00:00:40.48" resultid="7225" heatid="10571" lane="4" entrytime="00:00:40.20" entrycourse="LCM" />
                <RESULT eventid="1219" points="276" swimtime="00:01:27.33" resultid="7226" heatid="10593" lane="3" entrytime="00:01:29.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="187" swimtime="00:00:41.11" resultid="7227" heatid="10681" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Dominguez Olivieski" birthdate="2011-04-27" gender="M" nation="BRA" license="405717" swrid="5664737" athleteid="7243" externalid="405717">
              <RESULTS>
                <RESULT eventid="1103" points="295" swimtime="00:00:33.45" resultid="7244" heatid="10501" lane="9" />
                <RESULT eventid="1187" points="186" swimtime="00:00:45.45" resultid="7245" heatid="10571" lane="9" entrytime="00:00:44.87" entrycourse="LCM" />
                <RESULT eventid="1155" points="295" swimtime="00:01:09.63" resultid="7246" heatid="10540" lane="7" entrytime="00:01:13.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="318" swimtime="00:00:30.63" resultid="7247" heatid="10615" lane="9" entrytime="00:00:33.45" entrycourse="LCM" />
                <RESULT eventid="1219" points="185" swimtime="00:01:39.67" resultid="7248" heatid="10593" lane="9" entrytime="00:01:37.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="228" swimtime="00:00:38.54" resultid="7249" heatid="10684" lane="9" entrytime="00:00:42.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="14" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="AQUAFOZ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1203" points="250" swimtime="00:11:03.87" resultid="7257" heatid="10579" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                    <SPLIT distance="100" swimtime="00:01:09.15" />
                    <SPLIT distance="150" swimtime="00:01:49.31" />
                    <SPLIT distance="200" swimtime="00:02:29.99" />
                    <SPLIT distance="250" swimtime="00:03:09.48" />
                    <SPLIT distance="300" swimtime="00:03:54.24" />
                    <SPLIT distance="350" swimtime="00:04:40.07" />
                    <SPLIT distance="400" swimtime="00:05:23.42" />
                    <SPLIT distance="450" swimtime="00:05:59.99" />
                    <SPLIT distance="500" swimtime="00:06:42.25" />
                    <SPLIT distance="550" swimtime="00:07:31.02" />
                    <SPLIT distance="600" swimtime="00:08:18.97" />
                    <SPLIT distance="650" swimtime="00:08:54.00" />
                    <SPLIT distance="700" swimtime="00:09:34.30" />
                    <SPLIT distance="750" swimtime="00:10:19.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7228" number="1" />
                    <RELAYPOSITION athleteid="7223" number="2" />
                    <RELAYPOSITION athleteid="7233" number="3" />
                    <RELAYPOSITION athleteid="7238" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="AQUAFOZ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1325" points="263" swimtime="00:05:22.40" resultid="7258" heatid="10694" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.86" />
                    <SPLIT distance="150" swimtime="00:01:58.48" />
                    <SPLIT distance="200" swimtime="00:02:45.26" />
                    <SPLIT distance="250" swimtime="00:03:24.48" />
                    <SPLIT distance="300" swimtime="00:04:12.72" />
                    <SPLIT distance="350" swimtime="00:04:45.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7228" number="1" />
                    <RELAYPOSITION athleteid="7223" number="2" />
                    <RELAYPOSITION athleteid="7233" number="3" />
                    <RELAYPOSITION athleteid="7238" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1393" points="317" swimtime="00:04:35.79" resultid="7259" heatid="10750" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                    <SPLIT distance="100" swimtime="00:01:09.34" />
                    <SPLIT distance="150" swimtime="00:01:43.05" />
                    <SPLIT distance="200" swimtime="00:02:22.95" />
                    <SPLIT distance="250" swimtime="00:02:54.61" />
                    <SPLIT distance="300" swimtime="00:03:32.41" />
                    <SPLIT distance="350" swimtime="00:04:01.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7238" number="1" />
                    <RELAYPOSITION athleteid="7233" number="2" />
                    <RELAYPOSITION athleteid="7243" number="3" />
                    <RELAYPOSITION athleteid="7228" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="13025" nation="BRA" region="PR" clubid="7396" swrid="93779" name="Instituto Desportos Aquáticos De Foz Do Iguaçu" shortname="Cataratas Natação">
          <ATHLETES>
            <ATHLETE firstname="Bianca" lastname="Leticia Sbardelatti" birthdate="2011-07-28" gender="F" nation="BRA" license="403147" swrid="5676303" athleteid="7487" externalid="403147" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1179" points="256" swimtime="00:00:45.87" resultid="7488" heatid="10562" lane="0" entrytime="00:00:47.77" entrycourse="LCM" />
                <RESULT eventid="1147" points="337" swimtime="00:01:14.28" resultid="7489" heatid="10525" lane="6" entrytime="00:01:22.08" entrycourse="LCM" />
                <RESULT eventid="1227" points="360" swimtime="00:00:33.16" resultid="7490" heatid="10602" lane="8" entrytime="00:00:36.77" entrycourse="LCM" />
                <RESULT eventid="1297" points="229" swimtime="00:00:43.89" resultid="7491" heatid="10677" lane="5" entrytime="00:00:47.29" entrycourse="LCM" />
                <RESULT eventid="1281" points="245" swimtime="00:02:59.13" resultid="7492" heatid="10654" lane="7" entrytime="00:03:08.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.09" />
                    <SPLIT distance="100" swimtime="00:01:25.44" />
                    <SPLIT distance="150" swimtime="00:02:14.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Gabriel Dreher" birthdate="2011-12-05" gender="M" nation="BRA" license="403148" swrid="5676302" athleteid="7473" externalid="403148" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1187" points="173" swimtime="00:00:46.50" resultid="7474" heatid="10570" lane="3" entrytime="00:00:45.90" entrycourse="LCM" />
                <RESULT eventid="1155" points="276" swimtime="00:01:11.22" resultid="7475" heatid="10538" lane="2" entrytime="00:01:22.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="273" swimtime="00:00:32.23" resultid="7476" heatid="10614" lane="9" entrytime="00:00:35.68" entrycourse="LCM" />
                <RESULT eventid="1219" points="169" swimtime="00:01:42.83" resultid="7477" heatid="10590" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="270" swimtime="00:00:36.41" resultid="7478" heatid="10684" lane="7" entrytime="00:00:39.94" entrycourse="LCM" />
                <RESULT eventid="1289" points="280" swimtime="00:02:35.88" resultid="7479" heatid="10664" lane="5" entrytime="00:02:54.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.03" />
                    <SPLIT distance="100" swimtime="00:01:14.62" />
                    <SPLIT distance="150" swimtime="00:01:56.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Faisal" lastname="Basem Ghotme" birthdate="2010-12-18" gender="M" nation="BRA" license="390809" swrid="5596871" athleteid="7459" externalid="390809" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1071" points="421" swimtime="00:02:29.23" resultid="7460" heatid="10479" lane="8" entrytime="00:02:26.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                    <SPLIT distance="150" swimtime="00:01:50.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="489" swimtime="00:00:58.86" resultid="7461" heatid="10549" lane="1" entrytime="00:00:59.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="503" swimtime="00:00:26.28" resultid="7462" heatid="10625" lane="6" entrytime="00:00:26.17" entrycourse="LCM" />
                <RESULT eventid="1305" points="444" swimtime="00:00:30.85" resultid="7463" heatid="10686" lane="5" entrytime="00:00:30.58" entrycourse="LCM" />
                <RESULT eventid="1289" points="436" swimtime="00:02:14.45" resultid="7464" heatid="10669" lane="5" entrytime="00:02:19.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                    <SPLIT distance="100" swimtime="00:01:03.99" />
                    <SPLIT distance="150" swimtime="00:01:39.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="453" swimtime="00:01:07.17" resultid="7465" heatid="10740" lane="5" entrytime="00:01:06.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edward" lastname="Mikael De Lima" birthdate="2012-03-11" gender="M" nation="BRA" license="376445" swrid="5588816" athleteid="7507" externalid="376445" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1171" points="265" swimtime="00:02:51.76" resultid="7508" heatid="10555" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                    <SPLIT distance="100" swimtime="00:01:18.06" />
                    <SPLIT distance="150" swimtime="00:02:05.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="475" swimtime="00:00:59.46" resultid="7509" heatid="10546" lane="1" entrytime="00:01:02.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="454" swimtime="00:00:27.20" resultid="7510" heatid="10622" lane="5" entrytime="00:00:27.96" entrycourse="LCM" />
                <RESULT eventid="1289" points="461" swimtime="00:02:12.02" resultid="7511" heatid="10671" lane="1" entrytime="00:02:14.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.91" />
                    <SPLIT distance="100" swimtime="00:01:03.51" />
                    <SPLIT distance="150" swimtime="00:01:37.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="385" swimtime="00:01:07.96" resultid="7512" heatid="10706" lane="8" entrytime="00:01:19.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" status="DNS" swimtime="00:00:00.00" resultid="7513" heatid="10720" lane="7" entrytime="00:05:11.31" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanna" lastname="Mattiello" birthdate="2009-04-11" gender="F" nation="BRA" license="367011" swrid="5596914" athleteid="7445" externalid="367011" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1079" points="308" swimtime="00:03:23.56" resultid="7446" heatid="10481" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.38" />
                    <SPLIT distance="100" swimtime="00:01:37.29" />
                    <SPLIT distance="150" swimtime="00:02:31.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="357" swimtime="00:00:41.07" resultid="7447" heatid="10561" lane="6" />
                <RESULT eventid="1147" points="446" swimtime="00:01:07.68" resultid="7448" heatid="10530" lane="6" entrytime="00:01:08.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="450" swimtime="00:00:30.79" resultid="7449" heatid="10607" lane="8" entrytime="00:00:30.58" entrycourse="LCM" />
                <RESULT eventid="1281" points="432" swimtime="00:02:28.38" resultid="7450" heatid="10658" lane="8" entrytime="00:02:26.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                    <SPLIT distance="100" swimtime="00:01:12.10" />
                    <SPLIT distance="150" swimtime="00:01:51.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="400" swimtime="00:05:19.25" resultid="7451" heatid="10714" lane="8" entrytime="00:05:26.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                    <SPLIT distance="100" swimtime="00:01:18.64" />
                    <SPLIT distance="150" swimtime="00:02:01.16" />
                    <SPLIT distance="200" swimtime="00:02:41.55" />
                    <SPLIT distance="250" swimtime="00:03:22.00" />
                    <SPLIT distance="300" swimtime="00:04:01.96" />
                    <SPLIT distance="350" swimtime="00:04:42.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ysadora" lastname="Bertoldo" birthdate="2010-04-09" gender="F" nation="BRA" license="376444" swrid="5588553" athleteid="7493" externalid="376444" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1115" points="402" swimtime="00:20:46.30" resultid="7494" heatid="10511" lane="8" entrytime="00:20:10.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.98" />
                    <SPLIT distance="100" swimtime="00:01:15.28" />
                    <SPLIT distance="150" swimtime="00:01:56.06" />
                    <SPLIT distance="200" swimtime="00:02:36.75" />
                    <SPLIT distance="250" swimtime="00:03:18.34" />
                    <SPLIT distance="300" swimtime="00:03:59.41" />
                    <SPLIT distance="350" swimtime="00:04:40.67" />
                    <SPLIT distance="400" swimtime="00:05:21.97" />
                    <SPLIT distance="450" swimtime="00:06:04.07" />
                    <SPLIT distance="500" swimtime="00:06:46.16" />
                    <SPLIT distance="550" swimtime="00:07:28.03" />
                    <SPLIT distance="600" swimtime="00:08:10.11" />
                    <SPLIT distance="650" swimtime="00:08:52.52" />
                    <SPLIT distance="700" swimtime="00:09:34.35" />
                    <SPLIT distance="750" swimtime="00:10:16.31" />
                    <SPLIT distance="800" swimtime="00:10:58.53" />
                    <SPLIT distance="850" swimtime="00:11:40.92" />
                    <SPLIT distance="900" swimtime="00:12:23.48" />
                    <SPLIT distance="950" swimtime="00:13:05.47" />
                    <SPLIT distance="1000" swimtime="00:13:47.48" />
                    <SPLIT distance="1050" swimtime="00:14:30.20" />
                    <SPLIT distance="1100" swimtime="00:15:13.04" />
                    <SPLIT distance="1150" swimtime="00:15:55.92" />
                    <SPLIT distance="1200" swimtime="00:16:37.94" />
                    <SPLIT distance="1250" swimtime="00:17:20.49" />
                    <SPLIT distance="1300" swimtime="00:18:02.52" />
                    <SPLIT distance="1350" swimtime="00:18:44.66" />
                    <SPLIT distance="1400" swimtime="00:19:25.69" />
                    <SPLIT distance="1450" swimtime="00:20:06.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="352" swimtime="00:01:13.20" resultid="7495" heatid="10529" lane="2" entrytime="00:01:10.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="423" swimtime="00:10:45.60" resultid="7496" heatid="10632" lane="2" entrytime="00:10:33.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.60" />
                    <SPLIT distance="100" swimtime="00:01:15.13" />
                    <SPLIT distance="150" swimtime="00:01:55.09" />
                    <SPLIT distance="200" swimtime="00:02:36.42" />
                    <SPLIT distance="250" swimtime="00:03:17.25" />
                    <SPLIT distance="300" swimtime="00:03:58.41" />
                    <SPLIT distance="350" swimtime="00:04:39.41" />
                    <SPLIT distance="400" swimtime="00:05:20.53" />
                    <SPLIT distance="450" swimtime="00:06:01.94" />
                    <SPLIT distance="500" swimtime="00:06:43.22" />
                    <SPLIT distance="550" swimtime="00:07:24.30" />
                    <SPLIT distance="600" swimtime="00:08:05.92" />
                    <SPLIT distance="650" swimtime="00:08:46.67" />
                    <SPLIT distance="700" swimtime="00:09:27.35" />
                    <SPLIT distance="750" swimtime="00:10:07.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="389" swimtime="00:02:33.69" resultid="7497" heatid="10657" lane="6" entrytime="00:02:28.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                    <SPLIT distance="100" swimtime="00:01:15.70" />
                    <SPLIT distance="150" swimtime="00:01:55.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="409" swimtime="00:05:16.91" resultid="7498" heatid="10715" lane="8" entrytime="00:05:10.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                    <SPLIT distance="100" swimtime="00:01:15.14" />
                    <SPLIT distance="150" swimtime="00:01:55.64" />
                    <SPLIT distance="200" swimtime="00:02:36.69" />
                    <SPLIT distance="250" swimtime="00:03:17.65" />
                    <SPLIT distance="300" swimtime="00:03:58.25" />
                    <SPLIT distance="350" swimtime="00:04:38.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" status="DNS" swimtime="00:00:00.00" resultid="7499" heatid="10725" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Christopher" lastname="De Araujo" birthdate="2008-08-09" gender="M" nation="BRA" license="366376" swrid="5596884" athleteid="7431" externalid="366376" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1123" points="518" swimtime="00:09:22.61" resultid="7432" heatid="10513" lane="8" entrytime="00:09:13.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                    <SPLIT distance="100" swimtime="00:01:03.66" />
                    <SPLIT distance="150" swimtime="00:01:38.08" />
                    <SPLIT distance="200" swimtime="00:02:12.05" />
                    <SPLIT distance="250" swimtime="00:02:46.52" />
                    <SPLIT distance="300" swimtime="00:03:21.85" />
                    <SPLIT distance="350" swimtime="00:03:57.64" />
                    <SPLIT distance="400" swimtime="00:04:33.54" />
                    <SPLIT distance="450" swimtime="00:05:10.09" />
                    <SPLIT distance="500" swimtime="00:05:46.42" />
                    <SPLIT distance="550" swimtime="00:06:22.83" />
                    <SPLIT distance="600" swimtime="00:06:59.20" />
                    <SPLIT distance="650" swimtime="00:07:35.27" />
                    <SPLIT distance="700" swimtime="00:08:11.54" />
                    <SPLIT distance="750" swimtime="00:08:47.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="462" swimtime="00:05:13.65" resultid="7433" heatid="10522" lane="6" entrytime="00:05:19.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                    <SPLIT distance="100" swimtime="00:01:10.30" />
                    <SPLIT distance="150" swimtime="00:01:51.87" />
                    <SPLIT distance="200" swimtime="00:02:32.99" />
                    <SPLIT distance="250" swimtime="00:03:19.22" />
                    <SPLIT distance="300" swimtime="00:04:04.40" />
                    <SPLIT distance="350" swimtime="00:04:39.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" status="WDR" swimtime="00:00:00.00" resultid="7434" heatid="10635" lane="7" entrytime="00:17:44.18" entrycourse="LCM" />
                <RESULT eventid="1219" points="412" swimtime="00:01:16.44" resultid="7435" heatid="10598" lane="0" entrytime="00:01:13.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="491" swimtime="00:02:09.29" resultid="7436" heatid="10673" lane="2" entrytime="00:02:05.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.76" />
                    <SPLIT distance="100" swimtime="00:00:59.34" />
                    <SPLIT distance="150" swimtime="00:01:34.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="527" swimtime="00:04:32.44" resultid="7437" heatid="10723" lane="5" entrytime="00:04:28.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.57" />
                    <SPLIT distance="100" swimtime="00:01:00.57" />
                    <SPLIT distance="150" swimtime="00:01:35.01" />
                    <SPLIT distance="200" swimtime="00:02:10.30" />
                    <SPLIT distance="250" swimtime="00:02:46.34" />
                    <SPLIT distance="300" swimtime="00:03:22.47" />
                    <SPLIT distance="350" swimtime="00:03:58.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Axel" lastname="Ariel Giménez González" birthdate="2011-06-01" gender="M" nation="BRA" license="365755" swrid="5676299" athleteid="7452" externalid="365755" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1103" points="375" swimtime="00:00:30.88" resultid="7453" heatid="10499" lane="3" />
                <RESULT eventid="1187" points="348" swimtime="00:00:36.87" resultid="7454" heatid="10572" lane="6" entrytime="00:00:38.90" entrycourse="LCM" />
                <RESULT eventid="1155" points="431" swimtime="00:01:01.40" resultid="7455" heatid="10546" lane="7" entrytime="00:01:02.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="415" swimtime="00:00:28.02" resultid="7456" heatid="10621" lane="3" entrytime="00:00:28.51" entrycourse="LCM" />
                <RESULT eventid="1289" points="336" swimtime="00:02:26.61" resultid="7457" heatid="10666" lane="2" entrytime="00:02:35.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                    <SPLIT distance="100" swimtime="00:01:11.99" />
                    <SPLIT distance="150" swimtime="00:01:51.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="267" swimtime="00:01:20.08" resultid="7458" heatid="10736" lane="3" entrytime="00:01:20.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Marcio Peixoto" birthdate="2012-10-22" gender="M" nation="BRA" license="411994" swrid="5740013" athleteid="7500" externalid="411994">
              <RESULTS>
                <RESULT eventid="1103" points="145" swimtime="00:00:42.38" resultid="7501" heatid="10502" lane="9" />
                <RESULT eventid="1187" points="106" swimtime="00:00:54.67" resultid="7502" heatid="10569" lane="3" />
                <RESULT eventid="1155" points="231" swimtime="00:01:15.62" resultid="7503" heatid="10538" lane="6" entrytime="00:01:22.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="263" swimtime="00:00:32.60" resultid="7504" heatid="10613" lane="2" entrytime="00:00:38.65" entrycourse="LCM" />
                <RESULT eventid="1305" points="135" swimtime="00:00:45.88" resultid="7505" heatid="10683" lane="6" entrytime="00:00:52.23" entrycourse="LCM" />
                <RESULT eventid="1289" points="231" swimtime="00:02:46.23" resultid="7506" heatid="10664" lane="2" entrytime="00:03:01.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                    <SPLIT distance="150" swimtime="00:02:02.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Victor Oliveira" birthdate="2003-07-16" gender="M" nation="BRA" license="295723" swrid="5596944" athleteid="7417" externalid="295723" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1103" points="526" swimtime="00:00:27.58" resultid="7418" heatid="10508" lane="8" entrytime="00:00:27.54" entrycourse="LCM" />
                <RESULT eventid="1071" points="433" swimtime="00:02:27.88" resultid="7419" heatid="10480" lane="0" entrytime="00:02:22.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.17" />
                    <SPLIT distance="100" swimtime="00:01:11.19" />
                    <SPLIT distance="150" swimtime="00:01:49.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="351" swimtime="00:02:36.31" resultid="7420" heatid="10555" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                    <SPLIT distance="100" swimtime="00:01:04.66" />
                    <SPLIT distance="150" swimtime="00:01:44.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="487" swimtime="00:00:29.93" resultid="7421" heatid="10687" lane="2" entrytime="00:00:29.58" entrycourse="LCM" />
                <RESULT eventid="1341" points="486" swimtime="00:01:02.89" resultid="7422" heatid="10711" lane="9" entrytime="00:01:00.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="487" swimtime="00:01:05.56" resultid="7423" heatid="10742" lane="7" entrytime="00:01:03.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Monteiro Viebrantz" birthdate="2003-01-09" gender="M" nation="BRA" license="291175" swrid="5600219" athleteid="7407" externalid="291175">
              <RESULTS>
                <RESULT eventid="1235" points="615" swimtime="00:00:24.58" resultid="7408" heatid="10628" lane="9" entrytime="00:00:24.59" entrycourse="LCM" />
                <RESULT eventid="1305" points="501" swimtime="00:00:29.64" resultid="7409" heatid="10687" lane="8" entrytime="00:00:30.20" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Resende Ames" birthdate="2006-02-10" gender="M" nation="BRA" license="365657" swrid="5596931" athleteid="7424" externalid="365657" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1071" points="484" swimtime="00:02:22.45" resultid="7425" heatid="10479" lane="4" entrytime="00:02:24.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.71" />
                    <SPLIT distance="100" swimtime="00:01:09.93" />
                    <SPLIT distance="150" swimtime="00:01:46.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="499" swimtime="00:02:19.11" resultid="7426" heatid="10558" lane="5" entrytime="00:02:13.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.30" />
                    <SPLIT distance="100" swimtime="00:01:04.34" />
                    <SPLIT distance="150" swimtime="00:01:42.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="486" swimtime="00:05:08.37" resultid="7427" heatid="10522" lane="4" entrytime="00:05:13.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.30" />
                    <SPLIT distance="100" swimtime="00:01:03.50" />
                    <SPLIT distance="150" swimtime="00:01:42.41" />
                    <SPLIT distance="200" swimtime="00:02:22.13" />
                    <SPLIT distance="250" swimtime="00:03:12.65" />
                    <SPLIT distance="300" swimtime="00:04:01.88" />
                    <SPLIT distance="350" swimtime="00:04:34.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="509" swimtime="00:02:22.72" resultid="7428" heatid="10645" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.82" />
                    <SPLIT distance="100" swimtime="00:01:05.76" />
                    <SPLIT distance="150" swimtime="00:01:52.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="579" swimtime="00:00:59.30" resultid="7429" heatid="10711" lane="2" entrytime="00:00:59.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="478" swimtime="00:01:05.98" resultid="7430" heatid="10740" lane="1" entrytime="00:01:08.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Rogge" birthdate="2008-09-02" gender="M" nation="BRA" license="383387" swrid="4883279" athleteid="7410" externalid="383387" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1103" points="482" swimtime="00:00:28.40" resultid="7411" heatid="10506" lane="2" entrytime="00:00:30.40" entrycourse="LCM" />
                <RESULT eventid="1155" points="561" swimtime="00:00:56.24" resultid="7412" heatid="10550" lane="4" entrytime="00:00:56.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="552" swimtime="00:00:25.49" resultid="7413" heatid="10626" lane="5" entrytime="00:00:25.55" entrycourse="LCM" />
                <RESULT eventid="1305" points="398" swimtime="00:00:32.01" resultid="7414" heatid="10686" lane="1" entrytime="00:00:31.64" entrycourse="LCM" />
                <RESULT eventid="1289" points="377" swimtime="00:02:21.18" resultid="7415" heatid="10670" lane="3" entrytime="00:02:16.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                    <SPLIT distance="100" swimtime="00:01:08.21" />
                    <SPLIT distance="150" swimtime="00:01:45.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="343" swimtime="00:01:13.69" resultid="7416" heatid="10739" lane="9" entrytime="00:01:13.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Sermidi" birthdate="2005-06-15" gender="F" nation="BRA" license="283035" swrid="5596938" athleteid="7404" externalid="283035" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1227" points="450" swimtime="00:00:30.79" resultid="7405" heatid="10607" lane="6" entrytime="00:00:30.14" entrycourse="LCM" />
                <RESULT eventid="1297" points="369" swimtime="00:00:37.44" resultid="7406" heatid="10680" lane="9" entrytime="00:00:36.71" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Carvalho Carelli" birthdate="2011-10-15" gender="M" nation="BRA" license="403146" swrid="5676300" athleteid="7466" externalid="403146" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1103" points="407" swimtime="00:00:30.03" resultid="7467" heatid="10505" lane="5" entrytime="00:00:31.18" entrycourse="LCM" />
                <RESULT eventid="1171" points="346" swimtime="00:02:37.13" resultid="7468" heatid="10556" lane="9" entrytime="00:03:06.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                    <SPLIT distance="100" swimtime="00:01:12.45" />
                    <SPLIT distance="150" swimtime="00:01:55.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="382" swimtime="00:00:28.80" resultid="7469" heatid="10620" lane="7" entrytime="00:00:29.43" entrycourse="LCM" />
                <RESULT eventid="1289" points="461" swimtime="00:02:12.00" resultid="7470" heatid="10670" lane="9" entrytime="00:02:18.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.37" />
                    <SPLIT distance="100" swimtime="00:01:03.75" />
                    <SPLIT distance="150" swimtime="00:01:37.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="427" swimtime="00:01:05.62" resultid="7471" heatid="10707" lane="3" entrytime="00:01:12.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="358" swimtime="00:01:12.67" resultid="7472" heatid="10734" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Bailke" birthdate="2007-05-04" gender="M" nation="BRA" license="370566" swrid="5596869" athleteid="7438" externalid="370566" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1123" points="335" swimtime="00:10:50.85" resultid="7439" heatid="10515" lane="9" entrytime="00:10:34.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                    <SPLIT distance="100" swimtime="00:01:10.20" />
                    <SPLIT distance="150" swimtime="00:01:50.42" />
                    <SPLIT distance="200" swimtime="00:02:31.58" />
                    <SPLIT distance="250" swimtime="00:03:13.14" />
                    <SPLIT distance="300" swimtime="00:03:55.40" />
                    <SPLIT distance="350" swimtime="00:04:38.61" />
                    <SPLIT distance="400" swimtime="00:05:20.74" />
                    <SPLIT distance="450" swimtime="00:06:01.90" />
                    <SPLIT distance="500" swimtime="00:06:43.98" />
                    <SPLIT distance="550" swimtime="00:07:25.93" />
                    <SPLIT distance="600" swimtime="00:08:06.98" />
                    <SPLIT distance="650" swimtime="00:08:47.59" />
                    <SPLIT distance="700" swimtime="00:09:29.50" />
                    <SPLIT distance="750" swimtime="00:10:11.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="232" swimtime="00:02:59.46" resultid="7440" heatid="10556" lane="0" entrytime="00:03:03.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                    <SPLIT distance="100" swimtime="00:01:16.03" />
                    <SPLIT distance="150" swimtime="00:02:06.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="349" swimtime="00:20:35.86" resultid="7441" heatid="10637" lane="2" entrytime="00:20:31.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                    <SPLIT distance="100" swimtime="00:01:13.27" />
                    <SPLIT distance="150" swimtime="00:01:53.59" />
                    <SPLIT distance="200" swimtime="00:02:34.67" />
                    <SPLIT distance="250" swimtime="00:03:15.53" />
                    <SPLIT distance="300" swimtime="00:03:57.45" />
                    <SPLIT distance="350" swimtime="00:04:40.75" />
                    <SPLIT distance="400" swimtime="00:05:23.07" />
                    <SPLIT distance="450" swimtime="00:06:04.58" />
                    <SPLIT distance="500" swimtime="00:06:47.26" />
                    <SPLIT distance="550" swimtime="00:07:29.18" />
                    <SPLIT distance="600" swimtime="00:08:11.92" />
                    <SPLIT distance="650" swimtime="00:08:53.52" />
                    <SPLIT distance="700" swimtime="00:09:36.41" />
                    <SPLIT distance="750" swimtime="00:10:19.27" />
                    <SPLIT distance="800" swimtime="00:11:03.24" />
                    <SPLIT distance="850" swimtime="00:11:43.36" />
                    <SPLIT distance="900" swimtime="00:12:24.87" />
                    <SPLIT distance="950" swimtime="00:13:06.32" />
                    <SPLIT distance="1000" swimtime="00:13:46.83" />
                    <SPLIT distance="1050" swimtime="00:14:28.68" />
                    <SPLIT distance="1100" swimtime="00:15:11.32" />
                    <SPLIT distance="1150" swimtime="00:15:51.08" />
                    <SPLIT distance="1200" swimtime="00:16:32.47" />
                    <SPLIT distance="1250" swimtime="00:17:14.68" />
                    <SPLIT distance="1300" swimtime="00:17:56.61" />
                    <SPLIT distance="1350" swimtime="00:18:38.91" />
                    <SPLIT distance="1400" swimtime="00:19:21.45" />
                    <SPLIT distance="1450" swimtime="00:19:58.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="342" swimtime="00:00:29.88" resultid="7442" heatid="10613" lane="1" />
                <RESULT eventid="1341" points="340" swimtime="00:01:10.85" resultid="7443" heatid="10707" lane="4" entrytime="00:01:11.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="385" swimtime="00:05:02.34" resultid="7444" heatid="10720" lane="8" entrytime="00:05:12.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                    <SPLIT distance="100" swimtime="00:01:10.85" />
                    <SPLIT distance="150" swimtime="00:01:50.36" />
                    <SPLIT distance="200" swimtime="00:02:29.89" />
                    <SPLIT distance="250" swimtime="00:03:10.30" />
                    <SPLIT distance="300" swimtime="00:03:50.98" />
                    <SPLIT distance="350" swimtime="00:04:28.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Pinheiro" birthdate="2008-09-04" gender="F" nation="BRA" license="331610" swrid="5596894" athleteid="7397" externalid="331610">
              <RESULTS>
                <RESULT eventid="1063" points="404" swimtime="00:02:46.54" resultid="7398" heatid="10472" lane="6" entrytime="00:02:45.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.77" />
                    <SPLIT distance="100" swimtime="00:01:20.38" />
                    <SPLIT distance="150" swimtime="00:02:03.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="438" swimtime="00:05:48.12" resultid="7399" heatid="10520" lane="6" entrytime="00:05:47.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.84" />
                    <SPLIT distance="100" swimtime="00:01:16.81" />
                    <SPLIT distance="150" swimtime="00:02:01.55" />
                    <SPLIT distance="200" swimtime="00:02:45.32" />
                    <SPLIT distance="250" swimtime="00:03:38.41" />
                    <SPLIT distance="300" swimtime="00:04:30.21" />
                    <SPLIT distance="350" swimtime="00:05:10.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="430" swimtime="00:02:46.98" resultid="7400" heatid="10643" lane="1" entrytime="00:02:45.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                    <SPLIT distance="100" swimtime="00:01:18.17" />
                    <SPLIT distance="150" swimtime="00:02:10.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="422" swimtime="00:02:29.58" resultid="7401" heatid="10658" lane="7" entrytime="00:02:25.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                    <SPLIT distance="100" swimtime="00:01:12.62" />
                    <SPLIT distance="150" swimtime="00:01:51.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="397" swimtime="00:01:15.07" resultid="7402" heatid="10702" lane="8" entrytime="00:01:12.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="364" swimtime="00:01:20.00" resultid="7403" heatid="10731" lane="7" entrytime="00:01:16.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Resende Ames" birthdate="2010-02-02" gender="M" nation="BRA" license="365505" swrid="5588876" athleteid="7480" externalid="365505" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1071" points="450" swimtime="00:02:25.97" resultid="7481" heatid="10479" lane="2" entrytime="00:02:25.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                    <SPLIT distance="100" swimtime="00:01:10.98" />
                    <SPLIT distance="150" swimtime="00:01:48.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="400" swimtime="00:02:29.69" resultid="7482" heatid="10555" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="100" swimtime="00:01:09.77" />
                    <SPLIT distance="150" swimtime="00:01:50.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="396" swimtime="00:00:28.47" resultid="7483" heatid="10624" lane="6" entrytime="00:00:27.05" entrycourse="LCM" />
                <RESULT eventid="1305" points="417" swimtime="00:00:31.52" resultid="7484" heatid="10686" lane="2" entrytime="00:00:31.30" entrycourse="LCM" />
                <RESULT eventid="1341" points="410" swimtime="00:01:06.55" resultid="7485" heatid="10709" lane="8" entrytime="00:01:06.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="452" swimtime="00:01:07.20" resultid="7486" heatid="10740" lane="4" entrytime="00:01:06.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="19" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="CATARATAS &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1207" points="501" swimtime="00:08:46.72" resultid="7514" heatid="10581" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.84" />
                    <SPLIT distance="100" swimtime="00:00:58.82" />
                    <SPLIT distance="150" swimtime="00:01:31.27" />
                    <SPLIT distance="200" swimtime="00:02:04.33" />
                    <SPLIT distance="250" swimtime="00:02:34.14" />
                    <SPLIT distance="300" swimtime="00:03:07.69" />
                    <SPLIT distance="350" swimtime="00:03:40.66" />
                    <SPLIT distance="400" swimtime="00:04:13.29" />
                    <SPLIT distance="450" swimtime="00:04:42.62" />
                    <SPLIT distance="500" swimtime="00:05:16.92" />
                    <SPLIT distance="550" swimtime="00:05:54.35" />
                    <SPLIT distance="600" swimtime="00:06:30.24" />
                    <SPLIT distance="650" swimtime="00:07:01.09" />
                    <SPLIT distance="700" swimtime="00:07:35.53" />
                    <SPLIT distance="750" swimtime="00:08:10.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7431" number="1" />
                    <RELAYPOSITION athleteid="7424" number="2" />
                    <RELAYPOSITION athleteid="7410" number="3" />
                    <RELAYPOSITION athleteid="7438" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="CATARATAS &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1203" points="349" swimtime="00:09:54.45" resultid="7515" heatid="10579" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                    <SPLIT distance="100" swimtime="00:01:02.98" />
                    <SPLIT distance="150" swimtime="00:01:37.45" />
                    <SPLIT distance="200" swimtime="00:02:13.04" />
                    <SPLIT distance="250" swimtime="00:02:44.88" />
                    <SPLIT distance="300" swimtime="00:03:21.70" />
                    <SPLIT distance="350" swimtime="00:04:01.28" />
                    <SPLIT distance="400" swimtime="00:04:38.65" />
                    <SPLIT distance="450" swimtime="00:05:07.85" />
                    <SPLIT distance="500" swimtime="00:05:41.92" />
                    <SPLIT distance="550" swimtime="00:06:19.42" />
                    <SPLIT distance="600" swimtime="00:06:59.71" />
                    <SPLIT distance="650" swimtime="00:07:36.65" />
                    <SPLIT distance="700" swimtime="00:08:21.98" />
                    <SPLIT distance="750" swimtime="00:09:09.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7466" number="1" />
                    <RELAYPOSITION athleteid="7452" number="2" />
                    <RELAYPOSITION athleteid="7507" number="3" />
                    <RELAYPOSITION athleteid="7500" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="CATARATAS &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1331" points="511" swimtime="00:04:18.48" resultid="7516" heatid="10698" lane="6" entrytime="00:04:25.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="100" swimtime="00:01:06.06" />
                    <SPLIT distance="150" swimtime="00:01:42.24" />
                    <SPLIT distance="200" swimtime="00:02:22.77" />
                    <SPLIT distance="250" swimtime="00:02:51.23" />
                    <SPLIT distance="300" swimtime="00:03:21.51" />
                    <SPLIT distance="350" swimtime="00:03:48.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7417" number="1" />
                    <RELAYPOSITION athleteid="7431" number="2" />
                    <RELAYPOSITION athleteid="7424" number="3" />
                    <RELAYPOSITION athleteid="7410" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1399" points="565" swimtime="00:03:47.64" resultid="7518" heatid="10753" lane="2" entrytime="00:03:52.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.70" />
                    <SPLIT distance="100" swimtime="00:00:55.97" />
                    <SPLIT distance="150" swimtime="00:01:23.45" />
                    <SPLIT distance="200" swimtime="00:01:53.90" />
                    <SPLIT distance="250" swimtime="00:02:20.98" />
                    <SPLIT distance="300" swimtime="00:02:51.02" />
                    <SPLIT distance="350" swimtime="00:03:18.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7410" number="1" />
                    <RELAYPOSITION athleteid="7417" number="2" />
                    <RELAYPOSITION athleteid="7431" number="3" />
                    <RELAYPOSITION athleteid="7424" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="CATARATAS &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1325" points="366" swimtime="00:04:48.88" resultid="7517" heatid="10695" lane="2" entrytime="00:05:01.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                    <SPLIT distance="100" swimtime="00:01:19.65" />
                    <SPLIT distance="150" swimtime="00:01:57.16" />
                    <SPLIT distance="200" swimtime="00:02:41.33" />
                    <SPLIT distance="250" swimtime="00:03:12.52" />
                    <SPLIT distance="300" swimtime="00:03:48.56" />
                    <SPLIT distance="350" swimtime="00:04:16.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7473" number="1" />
                    <RELAYPOSITION athleteid="7452" number="2" />
                    <RELAYPOSITION athleteid="7466" number="3" />
                    <RELAYPOSITION athleteid="7507" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1393" points="385" swimtime="00:04:18.59" resultid="7519" heatid="10750" lane="2" entrytime="00:04:20.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                    <SPLIT distance="100" swimtime="00:01:03.33" />
                    <SPLIT distance="150" swimtime="00:01:32.92" />
                    <SPLIT distance="200" swimtime="00:02:05.25" />
                    <SPLIT distance="250" swimtime="00:02:33.38" />
                    <SPLIT distance="300" swimtime="00:03:03.95" />
                    <SPLIT distance="350" swimtime="00:03:39.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7452" number="1" />
                    <RELAYPOSITION athleteid="7466" number="2" />
                    <RELAYPOSITION athleteid="7507" number="3" />
                    <RELAYPOSITION athleteid="7500" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="X" name="CATARATAS &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1247" points="449" swimtime="00:04:43.78" resultid="7520" heatid="10631" lane="5" entrytime="00:04:30.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                    <SPLIT distance="100" swimtime="00:01:05.17" />
                    <SPLIT distance="150" swimtime="00:01:48.42" />
                    <SPLIT distance="200" swimtime="00:02:37.16" />
                    <SPLIT distance="250" swimtime="00:03:05.49" />
                    <SPLIT distance="300" swimtime="00:03:36.52" />
                    <SPLIT distance="350" swimtime="00:04:07.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7417" number="1" />
                    <RELAYPOSITION athleteid="7397" number="2" />
                    <RELAYPOSITION athleteid="7424" number="3" />
                    <RELAYPOSITION athleteid="7404" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="15969" nation="USA" clubid="8538" name="Estados Unidos da América" shortname="EUA">
          <ATHLETES>
            <ATHLETE firstname="Sophia" lastname="Alanis Whitney" birthdate="2007-07-21" gender="F" nation="USA" license="V397028" swrid="5757088" athleteid="8539" externalid="V397028">
              <RESULTS>
                <RESULT eventid="1095" points="509" status="EXH" swimtime="00:00:30.59" resultid="8540" heatid="10498" lane="3" entrytime="00:00:31.15" entrycourse="LCM" />
                <RESULT eventid="1147" points="487" status="EXH" swimtime="00:01:05.71" resultid="8541" heatid="10531" lane="2" entrytime="00:01:07.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="455" status="EXH" swimtime="00:00:30.68" resultid="8542" heatid="10607" lane="9" entrytime="00:00:30.62" entrycourse="LCM" />
                <RESULT eventid="1297" points="486" status="EXH" swimtime="00:00:34.16" resultid="8543" heatid="10680" lane="0" entrytime="00:00:35.70" entrycourse="LCM" />
                <RESULT eventid="1333" points="533" status="EXH" swimtime="00:01:08.02" resultid="8544" heatid="10702" lane="5" entrytime="00:01:07.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="453" status="EXH" swimtime="00:01:14.37" resultid="8545" heatid="10732" lane="1" entrytime="00:01:12.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="263" nation="BRA" region="PR" clubid="7820" swrid="75436" name="Clube Curitibano" shortname="Curitibano">
          <ATHLETES>
            <ATHLETE firstname="Rafael" lastname="Henrique Pasqual" birthdate="2005-05-07" gender="M" nation="BRA" license="329284" swrid="5600185" athleteid="8362" externalid="329284">
              <RESULTS>
                <RESULT eventid="1155" points="719" swimtime="00:00:51.79" resultid="8363" heatid="10552" lane="5" entrytime="00:00:52.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="680" swimtime="00:00:23.77" resultid="8364" heatid="10628" lane="5" entrytime="00:00:23.49" entrycourse="LCM" />
                <RESULT eventid="1289" points="632" swimtime="00:01:58.85" resultid="8365" heatid="10674" lane="1" entrytime="00:01:59.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.68" />
                    <SPLIT distance="100" swimtime="00:00:58.20" />
                    <SPLIT distance="150" swimtime="00:01:29.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Martynychen" birthdate="2011-12-19" gender="M" nation="BRA" license="366893" swrid="5602557" athleteid="8055" externalid="366893">
              <RESULTS>
                <RESULT eventid="1123" points="394" swimtime="00:10:16.49" resultid="8056" heatid="10514" lane="9" entrytime="00:10:02.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="100" swimtime="00:01:11.77" />
                    <SPLIT distance="150" swimtime="00:01:49.61" />
                    <SPLIT distance="200" swimtime="00:02:28.32" />
                    <SPLIT distance="250" swimtime="00:03:06.62" />
                    <SPLIT distance="300" swimtime="00:03:45.47" />
                    <SPLIT distance="350" swimtime="00:04:25.00" />
                    <SPLIT distance="400" swimtime="00:05:04.31" />
                    <SPLIT distance="450" swimtime="00:05:43.56" />
                    <SPLIT distance="500" swimtime="00:06:22.98" />
                    <SPLIT distance="550" swimtime="00:07:02.82" />
                    <SPLIT distance="600" swimtime="00:07:41.89" />
                    <SPLIT distance="650" swimtime="00:08:20.85" />
                    <SPLIT distance="700" swimtime="00:09:00.46" />
                    <SPLIT distance="750" swimtime="00:09:39.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="321" swimtime="00:02:43.32" resultid="8057" heatid="10477" lane="9" entrytime="00:02:45.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.96" />
                    <SPLIT distance="100" swimtime="00:01:18.46" />
                    <SPLIT distance="150" swimtime="00:02:01.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="301" swimtime="00:01:09.17" resultid="8058" heatid="10543" lane="2" entrytime="00:01:07.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="417" swimtime="00:19:24.68" resultid="8059" heatid="10636" lane="7" entrytime="00:19:12.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                    <SPLIT distance="100" swimtime="00:01:10.59" />
                    <SPLIT distance="150" swimtime="00:01:48.10" />
                    <SPLIT distance="200" swimtime="00:02:26.45" />
                    <SPLIT distance="250" swimtime="00:03:05.28" />
                    <SPLIT distance="300" swimtime="00:03:44.02" />
                    <SPLIT distance="350" swimtime="00:04:22.85" />
                    <SPLIT distance="400" swimtime="00:05:01.55" />
                    <SPLIT distance="450" swimtime="00:05:40.55" />
                    <SPLIT distance="500" swimtime="00:06:19.14" />
                    <SPLIT distance="550" swimtime="00:06:57.94" />
                    <SPLIT distance="600" swimtime="00:07:36.53" />
                    <SPLIT distance="650" swimtime="00:08:15.13" />
                    <SPLIT distance="700" swimtime="00:08:54.24" />
                    <SPLIT distance="750" swimtime="00:09:33.54" />
                    <SPLIT distance="800" swimtime="00:10:12.64" />
                    <SPLIT distance="850" swimtime="00:10:51.64" />
                    <SPLIT distance="900" swimtime="00:11:31.00" />
                    <SPLIT distance="950" swimtime="00:12:10.35" />
                    <SPLIT distance="1000" swimtime="00:12:49.88" />
                    <SPLIT distance="1050" swimtime="00:13:29.78" />
                    <SPLIT distance="1100" swimtime="00:14:09.24" />
                    <SPLIT distance="1150" swimtime="00:14:49.43" />
                    <SPLIT distance="1200" swimtime="00:15:28.34" />
                    <SPLIT distance="1250" swimtime="00:16:07.88" />
                    <SPLIT distance="1300" swimtime="00:16:47.18" />
                    <SPLIT distance="1350" swimtime="00:17:27.52" />
                    <SPLIT distance="1400" swimtime="00:18:06.80" />
                    <SPLIT distance="1450" swimtime="00:18:46.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="323" swimtime="00:02:28.57" resultid="8060" heatid="10668" lane="2" entrytime="00:02:22.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                    <SPLIT distance="100" swimtime="00:01:09.95" />
                    <SPLIT distance="150" swimtime="00:01:49.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="360" swimtime="00:05:09.17" resultid="8061" heatid="10721" lane="3" entrytime="00:04:53.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                    <SPLIT distance="100" swimtime="00:01:09.93" />
                    <SPLIT distance="150" swimtime="00:01:50.21" />
                    <SPLIT distance="200" swimtime="00:02:31.12" />
                    <SPLIT distance="250" swimtime="00:03:11.17" />
                    <SPLIT distance="300" swimtime="00:03:51.17" />
                    <SPLIT distance="350" swimtime="00:04:30.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Estevao" lastname="Valduga Artigas" birthdate="2009-06-01" gender="M" nation="BRA" license="339556" swrid="5600267" athleteid="7929" externalid="339556">
              <RESULTS>
                <RESULT eventid="1071" points="317" swimtime="00:02:44.08" resultid="7930" heatid="10476" lane="3" entrytime="00:02:46.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                    <SPLIT distance="100" swimtime="00:01:19.05" />
                    <SPLIT distance="150" swimtime="00:02:02.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="346" swimtime="00:00:29.76" resultid="7931" heatid="10618" lane="3" entrytime="00:00:30.48" entrycourse="LCM" />
                <RESULT eventid="1305" points="295" swimtime="00:00:35.35" resultid="7932" heatid="10684" lane="5" entrytime="00:00:37.08" entrycourse="LCM" />
                <RESULT eventid="1373" status="DNS" swimtime="00:00:00.00" resultid="7933" heatid="10737" lane="5" entrytime="00:01:16.31" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Valduga Artigas" birthdate="2009-06-01" gender="M" nation="BRA" license="339569" swrid="5600268" athleteid="7954" externalid="339569">
              <RESULTS>
                <RESULT eventid="1103" points="283" swimtime="00:00:33.91" resultid="7955" heatid="10505" lane="0" entrytime="00:00:32.57" entrycourse="LCM" />
                <RESULT eventid="1155" points="361" swimtime="00:01:05.14" resultid="7956" heatid="10544" lane="3" entrytime="00:01:06.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="360" swimtime="00:00:29.37" resultid="7957" heatid="10618" lane="6" entrytime="00:00:30.56" entrycourse="LCM" />
                <RESULT eventid="1341" status="DNS" swimtime="00:00:00.00" resultid="7958" heatid="10706" lane="6" entrytime="00:01:16.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Schiavon" birthdate="2010-05-03" gender="M" nation="BRA" license="356354" swrid="5600256" athleteid="8006" externalid="356354">
              <RESULTS>
                <RESULT eventid="1071" points="405" swimtime="00:02:31.18" resultid="8007" heatid="10478" lane="1" entrytime="00:02:31.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                    <SPLIT distance="100" swimtime="00:01:15.14" />
                    <SPLIT distance="150" swimtime="00:01:53.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="446" swimtime="00:05:17.27" resultid="8008" heatid="10522" lane="2" entrytime="00:05:19.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                    <SPLIT distance="100" swimtime="00:01:12.23" />
                    <SPLIT distance="150" swimtime="00:01:53.57" />
                    <SPLIT distance="200" swimtime="00:02:33.68" />
                    <SPLIT distance="250" swimtime="00:03:21.38" />
                    <SPLIT distance="300" swimtime="00:04:07.96" />
                    <SPLIT distance="350" swimtime="00:04:43.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="456" swimtime="00:02:28.08" resultid="8009" heatid="10650" lane="5" entrytime="00:02:30.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                    <SPLIT distance="100" swimtime="00:01:08.32" />
                    <SPLIT distance="150" swimtime="00:01:55.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="478" swimtime="00:02:10.38" resultid="8010" heatid="10671" lane="4" entrytime="00:02:10.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                    <SPLIT distance="100" swimtime="00:01:03.87" />
                    <SPLIT distance="150" swimtime="00:01:36.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="505" swimtime="00:04:36.28" resultid="8011" heatid="10723" lane="7" entrytime="00:04:35.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                    <SPLIT distance="100" swimtime="00:01:07.29" />
                    <SPLIT distance="150" swimtime="00:01:42.23" />
                    <SPLIT distance="200" swimtime="00:02:17.66" />
                    <SPLIT distance="250" swimtime="00:02:52.44" />
                    <SPLIT distance="300" swimtime="00:03:27.82" />
                    <SPLIT distance="350" swimtime="00:04:02.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="409" swimtime="00:01:09.49" resultid="8012" heatid="10739" lane="7" entrytime="00:01:11.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Coelho" birthdate="2011-11-11" gender="M" nation="BRA" license="366889" swrid="5602527" athleteid="8041" externalid="366889">
              <RESULTS>
                <RESULT eventid="1123" status="DNS" swimtime="00:00:00.00" resultid="8042" heatid="10515" lane="7" entrytime="00:10:22.54" entrycourse="LCM" />
                <RESULT eventid="1171" points="325" swimtime="00:02:40.35" resultid="8043" heatid="10556" lane="3" entrytime="00:02:43.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.87" />
                    <SPLIT distance="100" swimtime="00:01:16.24" />
                    <SPLIT distance="150" swimtime="00:01:59.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="433" swimtime="00:19:10.06" resultid="8044" heatid="10637" lane="6" entrytime="00:20:17.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                    <SPLIT distance="100" swimtime="00:01:13.91" />
                    <SPLIT distance="150" swimtime="00:01:52.53" />
                    <SPLIT distance="200" swimtime="00:02:30.81" />
                    <SPLIT distance="250" swimtime="00:03:08.97" />
                    <SPLIT distance="300" swimtime="00:03:47.34" />
                    <SPLIT distance="350" swimtime="00:04:26.08" />
                    <SPLIT distance="400" swimtime="00:05:04.53" />
                    <SPLIT distance="450" swimtime="00:05:42.89" />
                    <SPLIT distance="500" swimtime="00:06:21.23" />
                    <SPLIT distance="550" swimtime="00:07:00.16" />
                    <SPLIT distance="600" swimtime="00:07:38.47" />
                    <SPLIT distance="650" swimtime="00:08:17.27" />
                    <SPLIT distance="700" swimtime="00:08:56.14" />
                    <SPLIT distance="750" swimtime="00:09:34.64" />
                    <SPLIT distance="800" swimtime="00:10:13.27" />
                    <SPLIT distance="850" swimtime="00:10:52.60" />
                    <SPLIT distance="900" swimtime="00:11:31.32" />
                    <SPLIT distance="950" swimtime="00:12:10.05" />
                    <SPLIT distance="1000" swimtime="00:12:48.43" />
                    <SPLIT distance="1050" swimtime="00:13:27.33" />
                    <SPLIT distance="1100" swimtime="00:14:05.80" />
                    <SPLIT distance="1150" swimtime="00:14:44.21" />
                    <SPLIT distance="1200" swimtime="00:15:22.77" />
                    <SPLIT distance="1250" swimtime="00:16:01.52" />
                    <SPLIT distance="1300" swimtime="00:16:40.16" />
                    <SPLIT distance="1350" swimtime="00:17:19.10" />
                    <SPLIT distance="1400" swimtime="00:17:57.22" />
                    <SPLIT distance="1450" swimtime="00:18:35.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="420" swimtime="00:02:16.10" resultid="8045" heatid="10669" lane="6" entrytime="00:02:19.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                    <SPLIT distance="100" swimtime="00:01:06.64" />
                    <SPLIT distance="150" swimtime="00:01:42.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="338" swimtime="00:01:10.95" resultid="8046" heatid="10708" lane="8" entrytime="00:01:10.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="426" swimtime="00:04:52.41" resultid="8047" heatid="10721" lane="4" entrytime="00:04:53.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.43" />
                    <SPLIT distance="100" swimtime="00:01:08.75" />
                    <SPLIT distance="150" swimtime="00:01:46.45" />
                    <SPLIT distance="200" swimtime="00:02:24.33" />
                    <SPLIT distance="250" swimtime="00:03:02.23" />
                    <SPLIT distance="300" swimtime="00:03:40.27" />
                    <SPLIT distance="350" swimtime="00:04:17.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Prosdocimo" birthdate="2012-11-30" gender="M" nation="BRA" license="369272" swrid="5602575" athleteid="8182" externalid="369272">
              <RESULTS>
                <RESULT eventid="1123" points="335" swimtime="00:10:50.92" resultid="8183" heatid="10517" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.49" />
                    <SPLIT distance="100" swimtime="00:01:17.97" />
                    <SPLIT distance="200" swimtime="00:02:41.62" />
                    <SPLIT distance="250" swimtime="00:03:23.89" />
                    <SPLIT distance="300" swimtime="00:04:05.55" />
                    <SPLIT distance="350" swimtime="00:04:46.87" />
                    <SPLIT distance="400" swimtime="00:05:28.44" />
                    <SPLIT distance="450" swimtime="00:06:10.03" />
                    <SPLIT distance="500" swimtime="00:06:51.67" />
                    <SPLIT distance="550" swimtime="00:07:32.57" />
                    <SPLIT distance="600" swimtime="00:08:14.16" />
                    <SPLIT distance="650" swimtime="00:08:54.86" />
                    <SPLIT distance="700" swimtime="00:09:35.41" />
                    <SPLIT distance="750" swimtime="00:10:13.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="299" swimtime="00:02:47.31" resultid="8184" heatid="10476" lane="8" entrytime="00:02:52.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.58" />
                    <SPLIT distance="100" swimtime="00:01:22.27" />
                    <SPLIT distance="150" swimtime="00:02:06.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="307" swimtime="00:01:08.73" resultid="8185" heatid="10542" lane="4" entrytime="00:01:07.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="312" swimtime="00:00:30.80" resultid="8186" heatid="10616" lane="7" entrytime="00:00:32.06" entrycourse="LCM" />
                <RESULT eventid="1289" points="324" swimtime="00:02:28.38" resultid="8187" heatid="10667" lane="7" entrytime="00:02:29.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.46" />
                    <SPLIT distance="150" swimtime="00:01:51.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="314" swimtime="00:01:15.87" resultid="8188" heatid="10737" lane="9" entrytime="00:01:19.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Saboia" birthdate="2009-01-25" gender="M" nation="BRA" license="342252" swrid="5600253" athleteid="7944" externalid="342252">
              <RESULTS>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 10:53)" eventid="1087" status="DSQ" swimtime="00:02:41.71" resultid="7945" heatid="10492" lane="1" entrytime="00:02:38.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                    <SPLIT distance="100" swimtime="00:01:16.26" />
                    <SPLIT distance="150" swimtime="00:01:59.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="458" swimtime="00:00:33.66" resultid="7946" heatid="10574" lane="3" entrytime="00:00:33.69" entrycourse="LCM" />
                <RESULT eventid="1219" points="420" swimtime="00:01:15.95" resultid="7947" heatid="10598" lane="7" entrytime="00:01:12.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="424" swimtime="00:02:31.68" resultid="7948" heatid="10651" lane="9" entrytime="00:02:29.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                    <SPLIT distance="100" swimtime="00:01:13.87" />
                    <SPLIT distance="150" swimtime="00:01:57.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helen" lastname="Barato Bernardi" birthdate="2006-07-27" gender="F" nation="BRA" license="317031" swrid="5717244" athleteid="8349" externalid="317031">
              <RESULTS>
                <RESULT eventid="1079" points="650" swimtime="00:02:38.73" resultid="8350" heatid="10486" lane="4" entrytime="00:02:41.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.43" />
                    <SPLIT distance="100" swimtime="00:01:16.61" />
                    <SPLIT distance="150" swimtime="00:01:58.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nina" lastname="Rocha Ribeiro Da Silva" birthdate="2010-09-22" gender="F" nation="BRA" license="367216" swrid="5588884" athleteid="8298" externalid="367216">
              <RESULTS>
                <RESULT eventid="1079" points="430" swimtime="00:03:02.20" resultid="8299" heatid="10486" lane="9" entrytime="00:02:56.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.24" />
                    <SPLIT distance="100" swimtime="00:01:26.31" />
                    <SPLIT distance="150" swimtime="00:02:14.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="457" swimtime="00:00:37.84" resultid="8300" heatid="10565" lane="3" entrytime="00:00:35.76" entrycourse="LCM" />
                <RESULT eventid="1147" points="249" swimtime="00:01:22.13" resultid="8301" heatid="10531" lane="7" entrytime="00:01:07.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 9:45)" eventid="1227" status="DSQ" swimtime="00:00:38.12" resultid="8302" heatid="10606" lane="1" entrytime="00:00:31.06" entrycourse="LCM" />
                <RESULT eventid="1211" points="463" swimtime="00:01:22.85" resultid="8303" heatid="10589" lane="9" entrytime="00:01:20.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="380" swimtime="00:02:34.91" resultid="8304" heatid="10657" lane="7" entrytime="00:02:29.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                    <SPLIT distance="100" swimtime="00:01:14.67" />
                    <SPLIT distance="150" swimtime="00:01:54.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Bulla Lanaro" birthdate="2009-08-28" gender="F" nation="BRA" license="344301" swrid="5569976" athleteid="7865" externalid="344301">
              <RESULTS>
                <RESULT eventid="1095" points="549" swimtime="00:00:29.83" resultid="7866" heatid="10498" lane="4" entrytime="00:00:29.79" entrycourse="LCM" />
                <RESULT eventid="1163" points="507" swimtime="00:02:32.70" resultid="7867" heatid="10554" lane="4" entrytime="00:02:27.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                    <SPLIT distance="100" swimtime="00:01:10.83" />
                    <SPLIT distance="150" swimtime="00:01:52.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="583" swimtime="00:00:28.26" resultid="7868" heatid="10609" lane="5" entrytime="00:00:28.06" entrycourse="LCM" />
                <RESULT eventid="1281" points="590" swimtime="00:02:13.75" resultid="7869" heatid="10660" lane="5" entrytime="00:02:10.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.77" />
                    <SPLIT distance="100" swimtime="00:01:03.27" />
                    <SPLIT distance="150" swimtime="00:01:38.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="565" swimtime="00:01:06.74" resultid="7870" heatid="10702" lane="4" entrytime="00:01:04.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Xavier Jardim" birthdate="2012-01-23" gender="M" nation="BRA" license="369259" swrid="5641781" athleteid="8129" externalid="369259">
              <RESULTS>
                <RESULT eventid="1071" points="300" swimtime="00:02:47.17" resultid="8130" heatid="10476" lane="7" entrytime="00:02:50.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.06" />
                    <SPLIT distance="100" swimtime="00:01:21.28" />
                    <SPLIT distance="150" swimtime="00:02:05.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="352" swimtime="00:01:05.66" resultid="8131" heatid="10543" lane="9" entrytime="00:01:07.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="325" swimtime="00:00:30.39" resultid="8132" heatid="10617" lane="1" entrytime="00:00:31.34" entrycourse="LCM" />
                <RESULT eventid="1289" points="336" swimtime="00:02:26.58" resultid="8133" heatid="10666" lane="5" entrytime="00:02:34.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                    <SPLIT distance="100" swimtime="00:01:11.21" />
                    <SPLIT distance="150" swimtime="00:01:50.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="293" swimtime="00:01:17.68" resultid="8134" heatid="10737" lane="0" entrytime="00:01:19.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Brandt De Macedo" birthdate="2010-01-13" gender="M" nation="BRA" license="338925" swrid="5588565" athleteid="8027" externalid="338925">
              <RESULTS>
                <RESULT eventid="1123" points="513" swimtime="00:09:24.60" resultid="8028" heatid="10514" lane="5" entrytime="00:09:35.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                    <SPLIT distance="100" swimtime="00:01:06.62" />
                    <SPLIT distance="150" swimtime="00:01:41.72" />
                    <SPLIT distance="200" swimtime="00:02:17.28" />
                    <SPLIT distance="250" swimtime="00:02:52.80" />
                    <SPLIT distance="300" swimtime="00:03:28.33" />
                    <SPLIT distance="350" swimtime="00:04:04.19" />
                    <SPLIT distance="400" swimtime="00:04:40.20" />
                    <SPLIT distance="450" swimtime="00:05:15.75" />
                    <SPLIT distance="500" swimtime="00:05:51.76" />
                    <SPLIT distance="550" swimtime="00:06:27.80" />
                    <SPLIT distance="600" swimtime="00:07:03.66" />
                    <SPLIT distance="650" swimtime="00:07:39.93" />
                    <SPLIT distance="700" swimtime="00:08:15.74" />
                    <SPLIT distance="750" swimtime="00:08:51.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="452" swimtime="00:01:00.43" resultid="8029" heatid="10548" lane="4" entrytime="00:00:59.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="556" swimtime="00:17:38.73" resultid="8030" heatid="10635" lane="9" entrytime="00:18:34.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.31" />
                    <SPLIT distance="100" swimtime="00:01:05.67" />
                    <SPLIT distance="150" swimtime="00:01:40.26" />
                    <SPLIT distance="200" swimtime="00:02:15.49" />
                    <SPLIT distance="250" swimtime="00:02:50.68" />
                    <SPLIT distance="300" swimtime="00:03:25.97" />
                    <SPLIT distance="350" swimtime="00:04:01.34" />
                    <SPLIT distance="400" swimtime="00:04:37.10" />
                    <SPLIT distance="450" swimtime="00:05:12.60" />
                    <SPLIT distance="500" swimtime="00:05:47.97" />
                    <SPLIT distance="550" swimtime="00:06:23.33" />
                    <SPLIT distance="600" swimtime="00:06:59.01" />
                    <SPLIT distance="650" swimtime="00:07:34.67" />
                    <SPLIT distance="700" swimtime="00:08:10.39" />
                    <SPLIT distance="750" swimtime="00:08:45.81" />
                    <SPLIT distance="800" swimtime="00:09:21.55" />
                    <SPLIT distance="850" swimtime="00:09:56.98" />
                    <SPLIT distance="900" swimtime="00:10:32.72" />
                    <SPLIT distance="950" swimtime="00:11:08.39" />
                    <SPLIT distance="1000" swimtime="00:11:44.39" />
                    <SPLIT distance="1050" swimtime="00:12:19.91" />
                    <SPLIT distance="1100" swimtime="00:12:55.78" />
                    <SPLIT distance="1150" swimtime="00:13:31.21" />
                    <SPLIT distance="1200" swimtime="00:14:07.02" />
                    <SPLIT distance="1250" swimtime="00:14:42.56" />
                    <SPLIT distance="1300" swimtime="00:15:18.29" />
                    <SPLIT distance="1350" swimtime="00:15:53.99" />
                    <SPLIT distance="1400" swimtime="00:16:29.83" />
                    <SPLIT distance="1450" swimtime="00:17:04.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="398" swimtime="00:00:28.41" resultid="8031" heatid="10623" lane="2" entrytime="00:00:27.60" entrycourse="LCM" />
                <RESULT eventid="1289" points="444" swimtime="00:02:13.64" resultid="8032" heatid="10671" lane="3" entrytime="00:02:11.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.08" />
                    <SPLIT distance="100" swimtime="00:01:05.07" />
                    <SPLIT distance="150" swimtime="00:01:40.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="535" swimtime="00:04:31.07" resultid="8033" heatid="10723" lane="8" entrytime="00:04:37.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                    <SPLIT distance="100" swimtime="00:01:04.31" />
                    <SPLIT distance="150" swimtime="00:01:38.71" />
                    <SPLIT distance="200" swimtime="00:02:13.74" />
                    <SPLIT distance="250" swimtime="00:02:48.97" />
                    <SPLIT distance="300" swimtime="00:03:24.44" />
                    <SPLIT distance="350" swimtime="00:03:59.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Yolanda Ferreira" birthdate="2008-03-17" gender="F" nation="BRA" license="358335" swrid="5600276" athleteid="8249" externalid="358335">
              <RESULTS>
                <RESULT eventid="1079" points="503" swimtime="00:02:52.95" resultid="8250" heatid="10486" lane="2" entrytime="00:02:53.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                    <SPLIT distance="100" swimtime="00:01:22.97" />
                    <SPLIT distance="150" swimtime="00:02:08.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="508" swimtime="00:00:36.53" resultid="8251" heatid="10564" lane="5" entrytime="00:00:37.44" entrycourse="LCM" />
                <RESULT eventid="1227" points="493" swimtime="00:00:29.87" resultid="8252" heatid="10609" lane="0" entrytime="00:00:29.23" entrycourse="LCM" />
                <RESULT eventid="1211" points="482" swimtime="00:01:21.77" resultid="8253" heatid="10589" lane="1" entrytime="00:01:19.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="Pellanda" birthdate="2010-11-12" gender="M" nation="BRA" license="356352" swrid="5600233" athleteid="7913" externalid="356352">
              <RESULTS>
                <RESULT eventid="1123" status="DNS" swimtime="00:00:00.00" resultid="7914" heatid="10513" lane="5" entrytime="00:08:54.45" entrycourse="LCM" />
                <RESULT eventid="1155" status="DNS" swimtime="00:00:00.00" resultid="7915" heatid="10550" lane="2" entrytime="00:00:56.88" entrycourse="LCM" />
                <RESULT eventid="1257" status="DNS" swimtime="00:00:00.00" resultid="7916" heatid="10635" lane="4" entrytime="00:17:05.03" entrycourse="LCM" />
                <RESULT eventid="1235" status="DNS" swimtime="00:00:00.00" resultid="7917" heatid="10625" lane="7" entrytime="00:00:26.59" entrycourse="LCM" />
                <RESULT eventid="1289" status="DNS" swimtime="00:00:00.00" resultid="7918" heatid="10673" lane="3" entrytime="00:02:03.75" entrycourse="LCM" />
                <RESULT eventid="1357" status="DNS" swimtime="00:00:00.00" resultid="7919" heatid="10724" lane="2" entrytime="00:04:20.73" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabio" lastname="C Burak" birthdate="2009-08-29" gender="M" nation="BRA" license="343297" swrid="5600126" athleteid="8393" externalid="343297">
              <RESULTS>
                <RESULT eventid="1087" points="512" swimtime="00:02:36.83" resultid="8394" heatid="10492" lane="0" entrytime="00:02:39.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.73" />
                    <SPLIT distance="100" swimtime="00:01:16.43" />
                    <SPLIT distance="150" swimtime="00:01:57.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="504" swimtime="00:00:32.59" resultid="8395" heatid="10574" lane="4" entrytime="00:00:32.47" entrycourse="LCM" />
                <RESULT eventid="1219" points="510" swimtime="00:01:11.17" resultid="8396" heatid="10598" lane="2" entrytime="00:01:11.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="517" swimtime="00:02:21.97" resultid="8397" heatid="10652" lane="8" entrytime="00:02:21.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                    <SPLIT distance="100" swimtime="00:01:09.26" />
                    <SPLIT distance="150" swimtime="00:01:48.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="499" swimtime="00:01:05.05" resultid="8398" heatid="10741" lane="5" entrytime="00:01:04.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otavio" lastname="Araujo Barros" birthdate="2008-12-26" gender="M" nation="BRA" license="331713" swrid="5367497" athleteid="8118" externalid="331713">
              <RESULTS>
                <RESULT eventid="1123" points="595" swimtime="00:08:57.28" resultid="8119" heatid="10513" lane="6" entrytime="00:09:03.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.29" />
                    <SPLIT distance="100" swimtime="00:01:03.49" />
                    <SPLIT distance="150" swimtime="00:01:37.63" />
                    <SPLIT distance="200" swimtime="00:02:11.10" />
                    <SPLIT distance="250" swimtime="00:02:45.63" />
                    <SPLIT distance="300" swimtime="00:03:19.28" />
                    <SPLIT distance="350" swimtime="00:03:53.33" />
                    <SPLIT distance="400" swimtime="00:04:27.65" />
                    <SPLIT distance="450" swimtime="00:05:01.53" />
                    <SPLIT distance="500" swimtime="00:05:35.53" />
                    <SPLIT distance="550" swimtime="00:06:09.69" />
                    <SPLIT distance="600" swimtime="00:06:43.41" />
                    <SPLIT distance="650" swimtime="00:07:17.44" />
                    <SPLIT distance="700" swimtime="00:07:51.35" />
                    <SPLIT distance="750" swimtime="00:08:24.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="619" swimtime="00:01:59.62" resultid="8120" heatid="10674" lane="0" entrytime="00:02:00.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.13" />
                    <SPLIT distance="100" swimtime="00:00:58.72" />
                    <SPLIT distance="150" swimtime="00:01:29.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="619" swimtime="00:04:18.16" resultid="8121" heatid="10724" lane="3" entrytime="00:04:18.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                    <SPLIT distance="100" swimtime="00:01:01.70" />
                    <SPLIT distance="150" swimtime="00:01:34.17" />
                    <SPLIT distance="200" swimtime="00:02:06.83" />
                    <SPLIT distance="250" swimtime="00:02:39.71" />
                    <SPLIT distance="300" swimtime="00:03:12.47" />
                    <SPLIT distance="350" swimtime="00:03:46.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabelly" lastname="Sinnott" birthdate="2009-03-14" gender="F" nation="BRA" license="367255" swrid="5600258" athleteid="7859" externalid="367255">
              <RESULTS>
                <RESULT eventid="1115" points="593" swimtime="00:18:15.08" resultid="7860" heatid="10511" lane="6" entrytime="00:18:30.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                    <SPLIT distance="100" swimtime="00:01:08.82" />
                    <SPLIT distance="150" swimtime="00:01:44.79" />
                    <SPLIT distance="200" swimtime="00:02:20.60" />
                    <SPLIT distance="250" swimtime="00:02:56.83" />
                    <SPLIT distance="300" swimtime="00:03:33.04" />
                    <SPLIT distance="350" swimtime="00:04:09.81" />
                    <SPLIT distance="400" swimtime="00:04:46.23" />
                    <SPLIT distance="450" swimtime="00:05:22.78" />
                    <SPLIT distance="500" swimtime="00:05:59.34" />
                    <SPLIT distance="550" swimtime="00:06:35.78" />
                    <SPLIT distance="600" swimtime="00:07:12.27" />
                    <SPLIT distance="650" swimtime="00:07:48.85" />
                    <SPLIT distance="700" swimtime="00:08:25.43" />
                    <SPLIT distance="750" swimtime="00:09:01.95" />
                    <SPLIT distance="800" swimtime="00:09:38.44" />
                    <SPLIT distance="850" swimtime="00:10:15.10" />
                    <SPLIT distance="900" swimtime="00:10:51.68" />
                    <SPLIT distance="950" swimtime="00:11:28.52" />
                    <SPLIT distance="1000" swimtime="00:12:05.54" />
                    <SPLIT distance="1050" swimtime="00:12:42.62" />
                    <SPLIT distance="1100" swimtime="00:13:19.81" />
                    <SPLIT distance="1150" swimtime="00:13:57.19" />
                    <SPLIT distance="1200" swimtime="00:14:34.12" />
                    <SPLIT distance="1250" swimtime="00:15:11.14" />
                    <SPLIT distance="1300" swimtime="00:15:48.10" />
                    <SPLIT distance="1350" swimtime="00:16:25.21" />
                    <SPLIT distance="1400" swimtime="00:17:02.27" />
                    <SPLIT distance="1450" swimtime="00:17:39.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="626" swimtime="00:01:00.44" resultid="7861" heatid="10534" lane="3" entrytime="00:01:00.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="562" swimtime="00:09:47.11" resultid="7862" heatid="10632" lane="4" entrytime="00:09:50.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                    <SPLIT distance="100" swimtime="00:01:06.36" />
                    <SPLIT distance="150" swimtime="00:01:41.33" />
                    <SPLIT distance="200" swimtime="00:02:16.97" />
                    <SPLIT distance="250" swimtime="00:02:53.21" />
                    <SPLIT distance="300" swimtime="00:03:30.27" />
                    <SPLIT distance="350" swimtime="00:04:07.38" />
                    <SPLIT distance="400" swimtime="00:04:45.05" />
                    <SPLIT distance="450" swimtime="00:05:22.44" />
                    <SPLIT distance="500" swimtime="00:05:59.93" />
                    <SPLIT distance="550" swimtime="00:06:37.55" />
                    <SPLIT distance="600" swimtime="00:07:15.64" />
                    <SPLIT distance="650" swimtime="00:07:53.70" />
                    <SPLIT distance="700" swimtime="00:08:31.95" />
                    <SPLIT distance="750" swimtime="00:09:10.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="635" swimtime="00:02:10.53" resultid="7863" heatid="10660" lane="4" entrytime="00:02:09.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.93" />
                    <SPLIT distance="100" swimtime="00:01:02.30" />
                    <SPLIT distance="150" swimtime="00:01:35.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="605" swimtime="00:04:38.20" resultid="7864" heatid="10716" lane="4" entrytime="00:04:34.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                    <SPLIT distance="100" swimtime="00:01:07.76" />
                    <SPLIT distance="150" swimtime="00:01:41.95" />
                    <SPLIT distance="200" swimtime="00:02:16.17" />
                    <SPLIT distance="250" swimtime="00:02:50.89" />
                    <SPLIT distance="300" swimtime="00:03:26.36" />
                    <SPLIT distance="350" swimtime="00:04:02.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Fernandes" birthdate="2010-03-13" gender="M" nation="BRA" license="339266" swrid="5588695" athleteid="8307" externalid="339266">
              <RESULTS>
                <RESULT eventid="1071" points="401" swimtime="00:02:31.73" resultid="8308" heatid="10478" lane="3" entrytime="00:02:27.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                    <SPLIT distance="100" swimtime="00:01:11.20" />
                    <SPLIT distance="150" swimtime="00:01:50.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="518" swimtime="00:00:57.75" resultid="8309" heatid="10550" lane="8" entrytime="00:00:57.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="489" swimtime="00:00:26.54" resultid="8310" heatid="10625" lane="4" entrytime="00:00:26.09" entrycourse="LCM" />
                <RESULT eventid="1289" points="483" swimtime="00:02:09.99" resultid="8311" heatid="10673" lane="6" entrytime="00:02:04.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.66" />
                    <SPLIT distance="100" swimtime="00:01:01.35" />
                    <SPLIT distance="150" swimtime="00:01:35.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="452" swimtime="00:04:46.65" resultid="8312" heatid="10723" lane="0" entrytime="00:04:39.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.28" />
                    <SPLIT distance="100" swimtime="00:01:05.52" />
                    <SPLIT distance="150" swimtime="00:01:40.86" />
                    <SPLIT distance="200" swimtime="00:02:17.80" />
                    <SPLIT distance="250" swimtime="00:02:54.68" />
                    <SPLIT distance="300" swimtime="00:03:32.37" />
                    <SPLIT distance="350" swimtime="00:04:10.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="373" swimtime="00:01:11.66" resultid="8313" heatid="10740" lane="3" entrytime="00:01:07.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martina" lastname="Tallao Benke" birthdate="2012-01-02" gender="F" nation="BRA" license="376984" swrid="5588931" athleteid="8270" externalid="376984">
              <RESULTS>
                <RESULT eventid="1063" points="479" swimtime="00:02:37.29" resultid="8271" heatid="10473" lane="7" entrytime="00:02:37.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                    <SPLIT distance="100" swimtime="00:01:15.49" />
                    <SPLIT distance="150" swimtime="00:01:56.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="376" swimtime="00:02:48.70" resultid="8272" heatid="10554" lane="7" entrytime="00:02:53.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                    <SPLIT distance="100" swimtime="00:01:18.16" />
                    <SPLIT distance="150" swimtime="00:02:04.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="497" swimtime="00:00:29.80" resultid="8273" heatid="10608" lane="1" entrytime="00:00:29.64" entrycourse="LCM" />
                <RESULT eventid="1265" points="485" swimtime="00:02:40.51" resultid="8274" heatid="10643" lane="5" entrytime="00:02:43.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                    <SPLIT distance="100" swimtime="00:01:14.46" />
                    <SPLIT distance="150" swimtime="00:02:06.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="450" swimtime="00:01:12.00" resultid="8275" heatid="10702" lane="2" entrytime="00:01:11.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="476" swimtime="00:01:13.12" resultid="8276" heatid="10732" lane="3" entrytime="00:01:10.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carol" lastname="De Hertel" birthdate="2001-02-20" gender="F" nation="BRA" license="118424" swrid="5727648" athleteid="8360" externalid="118424">
              <RESULTS>
                <RESULT eventid="1115" points="594" swimtime="00:18:14.41" resultid="8361" heatid="10511" lane="4" entrytime="00:17:43.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.55" />
                    <SPLIT distance="100" swimtime="00:01:05.77" />
                    <SPLIT distance="150" swimtime="00:01:40.70" />
                    <SPLIT distance="200" swimtime="00:02:16.25" />
                    <SPLIT distance="250" swimtime="00:02:51.73" />
                    <SPLIT distance="300" swimtime="00:03:27.49" />
                    <SPLIT distance="350" swimtime="00:04:03.17" />
                    <SPLIT distance="400" swimtime="00:04:39.53" />
                    <SPLIT distance="450" swimtime="00:05:14.94" />
                    <SPLIT distance="500" swimtime="00:05:52.37" />
                    <SPLIT distance="550" swimtime="00:06:29.73" />
                    <SPLIT distance="600" swimtime="00:07:07.07" />
                    <SPLIT distance="650" swimtime="00:07:44.16" />
                    <SPLIT distance="700" swimtime="00:08:21.68" />
                    <SPLIT distance="750" swimtime="00:08:58.72" />
                    <SPLIT distance="800" swimtime="00:09:35.62" />
                    <SPLIT distance="850" swimtime="00:10:11.54" />
                    <SPLIT distance="900" swimtime="00:10:48.83" />
                    <SPLIT distance="950" swimtime="00:11:26.08" />
                    <SPLIT distance="1000" swimtime="00:12:03.55" />
                    <SPLIT distance="1050" swimtime="00:12:40.53" />
                    <SPLIT distance="1100" swimtime="00:13:17.63" />
                    <SPLIT distance="1150" swimtime="00:13:55.31" />
                    <SPLIT distance="1200" swimtime="00:14:32.50" />
                    <SPLIT distance="1250" swimtime="00:15:09.86" />
                    <SPLIT distance="1300" swimtime="00:15:47.04" />
                    <SPLIT distance="1350" swimtime="00:16:24.26" />
                    <SPLIT distance="1400" swimtime="00:17:01.30" />
                    <SPLIT distance="1450" swimtime="00:17:38.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Pereira Galle" birthdate="2011-08-02" gender="F" nation="BRA" license="369465" swrid="5627330" athleteid="8330" externalid="369465">
              <RESULTS>
                <RESULT eventid="1079" points="357" swimtime="00:03:13.77" resultid="8331" heatid="10484" lane="9" entrytime="00:03:07.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.54" />
                    <SPLIT distance="100" swimtime="00:01:32.62" />
                    <SPLIT distance="150" swimtime="00:02:23.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="361" swimtime="00:00:40.95" resultid="8332" heatid="10564" lane="6" entrytime="00:00:37.77" entrycourse="LCM" />
                <RESULT eventid="1147" points="409" swimtime="00:01:09.61" resultid="8333" heatid="10532" lane="9" entrytime="00:01:06.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="402" swimtime="00:00:31.97" resultid="8334" heatid="10606" lane="4" entrytime="00:00:30.69" entrycourse="LCM" />
                <RESULT eventid="1211" points="388" swimtime="00:01:27.86" resultid="8335" heatid="10588" lane="7" entrytime="00:01:22.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="409" swimtime="00:02:31.18" resultid="8336" heatid="10658" lane="9" entrytime="00:02:26.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                    <SPLIT distance="100" swimtime="00:01:13.06" />
                    <SPLIT distance="150" swimtime="00:01:52.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Clivatti" birthdate="2010-05-24" gender="M" nation="BRA" license="368007" swrid="5600139" athleteid="7901" externalid="368007">
              <RESULTS>
                <RESULT eventid="1123" points="519" swimtime="00:09:22.59" resultid="7902" heatid="10513" lane="9" entrytime="00:09:20.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.73" />
                    <SPLIT distance="100" swimtime="00:01:03.39" />
                    <SPLIT distance="150" swimtime="00:01:38.04" />
                    <SPLIT distance="200" swimtime="00:02:12.98" />
                    <SPLIT distance="250" swimtime="00:02:48.07" />
                    <SPLIT distance="300" swimtime="00:03:23.57" />
                    <SPLIT distance="350" swimtime="00:03:59.64" />
                    <SPLIT distance="400" swimtime="00:04:35.91" />
                    <SPLIT distance="450" swimtime="00:05:12.52" />
                    <SPLIT distance="500" swimtime="00:05:49.24" />
                    <SPLIT distance="550" swimtime="00:06:25.64" />
                    <SPLIT distance="600" swimtime="00:07:01.85" />
                    <SPLIT distance="650" swimtime="00:07:38.21" />
                    <SPLIT distance="700" swimtime="00:08:14.08" />
                    <SPLIT distance="750" swimtime="00:08:49.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="551" swimtime="00:00:56.57" resultid="7903" heatid="10550" lane="5" entrytime="00:00:56.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="504" swimtime="00:00:26.26" resultid="7904" heatid="10625" lane="2" entrytime="00:00:26.27" entrycourse="LCM" />
                <RESULT eventid="1289" points="571" swimtime="00:02:02.88" resultid="7905" heatid="10673" lane="5" entrytime="00:02:02.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.71" />
                    <SPLIT distance="100" swimtime="00:00:58.28" />
                    <SPLIT distance="150" swimtime="00:01:30.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="557" swimtime="00:04:27.35" resultid="7906" heatid="10724" lane="0" entrytime="00:04:25.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.44" />
                    <SPLIT distance="100" swimtime="00:01:02.89" />
                    <SPLIT distance="150" swimtime="00:01:36.86" />
                    <SPLIT distance="200" swimtime="00:02:10.98" />
                    <SPLIT distance="250" swimtime="00:02:45.73" />
                    <SPLIT distance="300" swimtime="00:03:20.31" />
                    <SPLIT distance="350" swimtime="00:03:54.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="278" swimtime="00:01:18.99" resultid="7907" heatid="10739" lane="0" entrytime="00:01:12.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Peret Saboia" birthdate="2009-11-25" gender="F" nation="BRA" license="342238" swrid="5600234" athleteid="7934" externalid="342238">
              <RESULTS>
                <RESULT eventid="1079" points="493" swimtime="00:02:54.11" resultid="7935" heatid="10486" lane="7" entrytime="00:02:54.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.10" />
                    <SPLIT distance="100" swimtime="00:01:23.47" />
                    <SPLIT distance="150" swimtime="00:02:09.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="465" swimtime="00:00:37.62" resultid="7936" heatid="10564" lane="4" entrytime="00:00:37.40" entrycourse="LCM" />
                <RESULT eventid="1211" points="509" swimtime="00:01:20.28" resultid="7937" heatid="10589" lane="6" entrytime="00:01:18.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="388" swimtime="00:01:18.30" resultid="7938" heatid="10725" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Rocha Silva" birthdate="2007-10-10" gender="M" nation="BRA" license="372280" swrid="5717294" athleteid="7889" externalid="372280">
              <RESULTS>
                <RESULT eventid="1155" points="759" swimtime="00:00:50.86" resultid="7890" heatid="10552" lane="4" entrytime="00:00:49.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="676" swimtime="00:00:23.82" resultid="7891" heatid="10628" lane="4" entrytime="00:00:23.39" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Emili Gomes Xavier" birthdate="2010-09-08" gender="F" nation="BRA" license="372519" swrid="5717260" athleteid="7922" externalid="372519">
              <RESULTS>
                <RESULT eventid="1095" points="282" swimtime="00:00:37.25" resultid="7923" heatid="10493" lane="6" />
                <RESULT eventid="1179" points="424" swimtime="00:00:38.81" resultid="7924" heatid="10561" lane="5" />
                <RESULT eventid="1147" points="528" swimtime="00:01:03.97" resultid="7925" heatid="10534" lane="8" entrytime="00:01:03.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="471" swimtime="00:00:30.33" resultid="7926" heatid="10608" lane="3" entrytime="00:00:29.33" entrycourse="LCM" />
                <RESULT eventid="1281" points="535" swimtime="00:02:18.23" resultid="7927" heatid="10659" lane="4" entrytime="00:02:20.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.76" />
                    <SPLIT distance="100" swimtime="00:01:06.44" />
                    <SPLIT distance="150" swimtime="00:01:43.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="501" swimtime="00:04:56.19" resultid="7928" heatid="10715" lane="7" entrytime="00:05:06.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                    <SPLIT distance="100" swimtime="00:01:10.20" />
                    <SPLIT distance="150" swimtime="00:01:48.48" />
                    <SPLIT distance="200" swimtime="00:02:25.97" />
                    <SPLIT distance="250" swimtime="00:03:04.14" />
                    <SPLIT distance="300" swimtime="00:03:42.11" />
                    <SPLIT distance="350" swimtime="00:04:20.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Albuquerque" birthdate="2012-11-16" gender="F" nation="BRA" license="369281" swrid="5602506" athleteid="8221" externalid="369281">
              <RESULTS>
                <RESULT eventid="1115" points="415" swimtime="00:20:33.84" resultid="8222" heatid="10512" lane="1" entrytime="00:21:44.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                    <SPLIT distance="100" swimtime="00:01:15.89" />
                    <SPLIT distance="150" swimtime="00:01:56.71" />
                    <SPLIT distance="200" swimtime="00:02:37.92" />
                    <SPLIT distance="250" swimtime="00:03:18.78" />
                    <SPLIT distance="300" swimtime="00:04:00.09" />
                    <SPLIT distance="350" swimtime="00:04:41.43" />
                    <SPLIT distance="400" swimtime="00:05:23.33" />
                    <SPLIT distance="450" swimtime="00:06:05.01" />
                    <SPLIT distance="500" swimtime="00:06:46.55" />
                    <SPLIT distance="550" swimtime="00:07:28.72" />
                    <SPLIT distance="600" swimtime="00:08:10.46" />
                    <SPLIT distance="650" swimtime="00:08:52.01" />
                    <SPLIT distance="700" swimtime="00:09:33.81" />
                    <SPLIT distance="750" swimtime="00:10:15.01" />
                    <SPLIT distance="800" swimtime="00:10:56.70" />
                    <SPLIT distance="850" swimtime="00:11:38.22" />
                    <SPLIT distance="900" swimtime="00:12:20.50" />
                    <SPLIT distance="950" swimtime="00:13:02.38" />
                    <SPLIT distance="1000" swimtime="00:13:43.97" />
                    <SPLIT distance="1050" swimtime="00:14:25.94" />
                    <SPLIT distance="1100" swimtime="00:15:07.83" />
                    <SPLIT distance="1150" swimtime="00:15:50.05" />
                    <SPLIT distance="1200" swimtime="00:16:31.68" />
                    <SPLIT distance="1250" swimtime="00:17:13.37" />
                    <SPLIT distance="1300" swimtime="00:17:55.25" />
                    <SPLIT distance="1350" swimtime="00:18:36.41" />
                    <SPLIT distance="1400" swimtime="00:19:17.29" />
                    <SPLIT distance="1450" swimtime="00:19:56.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="398" swimtime="00:03:06.89" resultid="8223" heatid="10483" lane="1" entrytime="00:03:16.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.08" />
                    <SPLIT distance="100" swimtime="00:01:31.00" />
                    <SPLIT distance="150" swimtime="00:02:19.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="401" swimtime="00:05:58.49" resultid="8224" heatid="10520" lane="8" entrytime="00:06:00.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                    <SPLIT distance="100" swimtime="00:01:25.82" />
                    <SPLIT distance="150" swimtime="00:02:14.36" />
                    <SPLIT distance="200" swimtime="00:03:00.77" />
                    <SPLIT distance="250" swimtime="00:03:51.04" />
                    <SPLIT distance="300" swimtime="00:04:40.21" />
                    <SPLIT distance="350" swimtime="00:05:20.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="409" swimtime="00:10:52.80" resultid="8225" heatid="10633" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.31" />
                    <SPLIT distance="100" swimtime="00:01:15.51" />
                    <SPLIT distance="150" swimtime="00:01:56.95" />
                    <SPLIT distance="200" swimtime="00:02:38.50" />
                    <SPLIT distance="250" swimtime="00:03:19.82" />
                    <SPLIT distance="300" swimtime="00:04:01.34" />
                    <SPLIT distance="350" swimtime="00:04:43.44" />
                    <SPLIT distance="400" swimtime="00:05:25.30" />
                    <SPLIT distance="450" swimtime="00:06:06.87" />
                    <SPLIT distance="500" swimtime="00:06:48.76" />
                    <SPLIT distance="550" swimtime="00:07:30.54" />
                    <SPLIT distance="600" swimtime="00:08:12.22" />
                    <SPLIT distance="650" swimtime="00:08:53.58" />
                    <SPLIT distance="700" swimtime="00:09:35.60" />
                    <SPLIT distance="750" swimtime="00:10:14.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="376" swimtime="00:01:28.80" resultid="8226" heatid="10586" lane="8" entrytime="00:01:30.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="394" swimtime="00:02:51.93" resultid="8227" heatid="10641" lane="5" entrytime="00:02:55.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.14" />
                    <SPLIT distance="100" swimtime="00:01:25.07" />
                    <SPLIT distance="150" swimtime="00:02:14.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Braun Prado" birthdate="2008-04-07" gender="M" nation="BRA" license="307663" swrid="5484324" athleteid="7965" externalid="307663">
              <RESULTS>
                <RESULT eventid="1071" points="512" swimtime="00:02:19.81" resultid="7966" heatid="10480" lane="3" entrytime="00:02:14.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                    <SPLIT distance="100" swimtime="00:01:07.75" />
                    <SPLIT distance="150" swimtime="00:01:43.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="497" swimtime="00:02:23.91" resultid="7967" heatid="10651" lane="1" entrytime="00:02:27.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.04" />
                    <SPLIT distance="100" swimtime="00:01:07.02" />
                    <SPLIT distance="150" swimtime="00:01:50.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="550" swimtime="00:01:02.96" resultid="7968" heatid="10742" lane="6" entrytime="00:01:01.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolau" lastname="Neto" birthdate="2011-03-22" gender="M" nation="BRA" license="366906" swrid="5602565" athleteid="8090" externalid="366906">
              <RESULTS>
                <RESULT eventid="1087" points="392" swimtime="00:02:51.43" resultid="8091" heatid="10490" lane="4" entrytime="00:02:53.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                    <SPLIT distance="100" swimtime="00:01:19.99" />
                    <SPLIT distance="150" swimtime="00:02:05.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="396" swimtime="00:00:35.32" resultid="8092" heatid="10573" lane="3" entrytime="00:00:35.75" entrycourse="LCM" />
                <RESULT eventid="1155" points="454" swimtime="00:01:00.37" resultid="8093" heatid="10547" lane="5" entrytime="00:01:01.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="435" swimtime="00:00:27.59" resultid="8094" heatid="10623" lane="9" entrytime="00:00:27.86" entrycourse="LCM" />
                <RESULT eventid="1219" points="416" swimtime="00:01:16.14" resultid="8095" heatid="10596" lane="5" entrytime="00:01:18.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="425" swimtime="00:02:15.61" resultid="8096" heatid="10669" lane="3" entrytime="00:02:19.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                    <SPLIT distance="100" swimtime="00:01:05.31" />
                    <SPLIT distance="150" swimtime="00:01:40.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Estela" lastname="Albuquerque" birthdate="2010-11-23" gender="F" nation="BRA" license="356344" swrid="5653285" athleteid="7992" externalid="356344">
              <RESULTS>
                <RESULT eventid="1147" points="427" swimtime="00:01:08.62" resultid="7993" heatid="10532" lane="1" entrytime="00:01:06.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="433" swimtime="00:00:31.19" resultid="7994" heatid="10605" lane="5" entrytime="00:00:31.26" entrycourse="LCM" />
                <RESULT eventid="1265" points="402" swimtime="00:02:50.87" resultid="7995" heatid="10641" lane="6" entrytime="00:02:59.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                    <SPLIT distance="100" swimtime="00:01:20.57" />
                    <SPLIT distance="150" swimtime="00:02:14.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="430" swimtime="00:02:28.66" resultid="7996" heatid="10659" lane="5" entrytime="00:02:21.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                    <SPLIT distance="100" swimtime="00:01:10.99" />
                    <SPLIT distance="150" swimtime="00:01:50.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="419" swimtime="00:05:14.52" resultid="7997" heatid="10716" lane="7" entrytime="00:04:58.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                    <SPLIT distance="100" swimtime="00:01:13.85" />
                    <SPLIT distance="150" swimtime="00:01:53.26" />
                    <SPLIT distance="200" swimtime="00:02:33.30" />
                    <SPLIT distance="250" swimtime="00:03:13.74" />
                    <SPLIT distance="300" swimtime="00:03:54.52" />
                    <SPLIT distance="350" swimtime="00:04:35.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="350" swimtime="00:01:21.06" resultid="7998" heatid="10730" lane="6" entrytime="00:01:18.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="De Czarnecki" birthdate="2008-06-24" gender="M" nation="BRA" license="329641" swrid="5600146" athleteid="7835" externalid="329641">
              <RESULTS>
                <RESULT eventid="1071" status="DNS" swimtime="00:00:00.00" resultid="7836" heatid="10480" lane="4" entrytime="00:02:11.87" entrycourse="LCM" />
                <RESULT eventid="1155" status="DNS" swimtime="00:00:00.00" resultid="7837" heatid="10552" lane="7" entrytime="00:00:53.65" entrycourse="LCM" />
                <RESULT eventid="1289" status="DNS" swimtime="00:00:00.00" resultid="7838" heatid="10674" lane="7" entrytime="00:01:58.81" entrycourse="LCM" />
                <RESULT eventid="1373" status="DNS" swimtime="00:00:00.00" resultid="7839" heatid="10742" lane="3" entrytime="00:01:00.97" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ricardo" lastname="De Lima Cavalcanti" birthdate="2009-12-17" gender="M" nation="BRA" license="380965" swrid="5634589" athleteid="8344" externalid="380965">
              <RESULTS>
                <RESULT eventid="1103" points="550" swimtime="00:00:27.17" resultid="8345" heatid="10508" lane="7" entrytime="00:00:27.23" entrycourse="LCM" />
                <RESULT eventid="1171" points="430" swimtime="00:02:26.15" resultid="8346" heatid="10558" lane="2" entrytime="00:02:21.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.59" />
                    <SPLIT distance="100" swimtime="00:01:06.48" />
                    <SPLIT distance="150" swimtime="00:01:45.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="501" swimtime="00:00:26.32" resultid="8347" heatid="10627" lane="6" entrytime="00:00:25.20" entrycourse="LCM" />
                <RESULT eventid="1341" points="509" swimtime="00:01:01.91" resultid="8348" heatid="10711" lane="8" entrytime="00:00:59.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Fernando Deschamps" birthdate="2006-01-20" gender="M" nation="BRA" license="352911" swrid="5811243" athleteid="8390" externalid="352911">
              <RESULTS>
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="8391" heatid="10575" lane="3" entrytime="00:00:29.39" entrycourse="LCM" />
                <RESULT eventid="1219" status="DNS" swimtime="00:00:00.00" resultid="8392" heatid="10599" lane="5" entrytime="00:01:04.08" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="De Almeida Dias" birthdate="2012-02-18" gender="F" nation="BRA" license="369262" swrid="5588638" athleteid="8142" externalid="369262">
              <RESULTS>
                <RESULT eventid="1063" points="351" swimtime="00:02:54.43" resultid="8143" heatid="10471" lane="7" entrytime="00:02:53.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.95" />
                    <SPLIT distance="100" swimtime="00:01:25.60" />
                    <SPLIT distance="150" swimtime="00:02:11.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="527" swimtime="00:01:03.99" resultid="8144" heatid="10532" lane="6" entrytime="00:01:05.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="405" swimtime="00:10:54.91" resultid="8145" heatid="10634" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                    <SPLIT distance="100" swimtime="00:01:15.97" />
                    <SPLIT distance="150" swimtime="00:01:57.38" />
                    <SPLIT distance="200" swimtime="00:02:39.80" />
                    <SPLIT distance="250" swimtime="00:03:21.21" />
                    <SPLIT distance="300" swimtime="00:04:03.26" />
                    <SPLIT distance="350" swimtime="00:04:45.24" />
                    <SPLIT distance="400" swimtime="00:05:26.57" />
                    <SPLIT distance="450" swimtime="00:06:08.55" />
                    <SPLIT distance="500" swimtime="00:06:50.17" />
                    <SPLIT distance="550" swimtime="00:07:31.74" />
                    <SPLIT distance="600" swimtime="00:08:13.79" />
                    <SPLIT distance="650" swimtime="00:08:55.08" />
                    <SPLIT distance="700" swimtime="00:09:36.43" />
                    <SPLIT distance="750" swimtime="00:10:16.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="385" swimtime="00:01:28.10" resultid="8146" heatid="10586" lane="1" entrytime="00:01:29.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="506" swimtime="00:02:20.83" resultid="8147" heatid="10659" lane="7" entrytime="00:02:22.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                    <SPLIT distance="100" swimtime="00:01:08.36" />
                    <SPLIT distance="150" swimtime="00:01:45.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="455" swimtime="00:05:05.97" resultid="8148" heatid="10715" lane="4" entrytime="00:05:03.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="100" swimtime="00:01:12.29" />
                    <SPLIT distance="150" swimtime="00:01:51.49" />
                    <SPLIT distance="200" swimtime="00:02:30.90" />
                    <SPLIT distance="250" swimtime="00:03:10.68" />
                    <SPLIT distance="300" swimtime="00:03:49.94" />
                    <SPLIT distance="350" swimtime="00:04:29.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Guimaraes E Souza" birthdate="2008-12-21" gender="M" nation="BRA" license="376972" swrid="5600182" athleteid="8266" externalid="376972">
              <RESULTS>
                <RESULT eventid="1087" points="542" swimtime="00:02:33.85" resultid="8267" heatid="10492" lane="7" entrytime="00:02:37.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                    <SPLIT distance="100" swimtime="00:01:15.45" />
                    <SPLIT distance="150" swimtime="00:01:55.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="581" swimtime="00:01:08.13" resultid="8268" heatid="10599" lane="0" entrytime="00:01:07.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="527" swimtime="00:02:21.12" resultid="8269" heatid="10651" lane="5" entrytime="00:02:24.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                    <SPLIT distance="100" swimtime="00:01:10.09" />
                    <SPLIT distance="150" swimtime="00:01:50.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Atihe Gomes" birthdate="2011-07-08" gender="F" nation="BRA" license="421515" swrid="5636897" athleteid="8401" externalid="421515">
              <RESULTS>
                <RESULT eventid="1179" points="198" swimtime="00:00:50.00" resultid="8402" heatid="10560" lane="3" />
                <RESULT eventid="1147" points="249" swimtime="00:01:22.15" resultid="8403" heatid="10526" lane="9" entrytime="00:01:20.92" entrycourse="LCM" />
                <RESULT eventid="1227" points="276" swimtime="00:00:36.22" resultid="8404" heatid="10602" lane="7" entrytime="00:00:35.58" entrycourse="LCM" />
                <RESULT eventid="1211" points="219" swimtime="00:01:46.38" resultid="8405" heatid="10583" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Fontolan Gomes" birthdate="2010-07-02" gender="M" nation="BRA" license="356245" swrid="5588705" athleteid="7978" externalid="356245">
              <RESULTS>
                <RESULT eventid="1071" points="380" swimtime="00:02:34.51" resultid="7979" heatid="10478" lane="7" entrytime="00:02:31.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="100" swimtime="00:01:13.88" />
                    <SPLIT distance="150" swimtime="00:01:54.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="343" swimtime="00:01:06.27" resultid="7980" heatid="10544" lane="7" entrytime="00:01:06.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" status="DNS" swimtime="00:00:00.00" resultid="7981" heatid="10616" lane="3" entrytime="00:00:31.96" entrycourse="LCM" />
                <RESULT eventid="1219" status="DNS" swimtime="00:00:00.00" resultid="7982" heatid="10593" lane="2" entrytime="00:01:31.02" entrycourse="LCM" />
                <RESULT eventid="1289" status="DNS" swimtime="00:00:00.00" resultid="7983" heatid="10669" lane="9" entrytime="00:02:20.23" entrycourse="LCM" />
                <RESULT eventid="1373" status="DNS" swimtime="00:00:00.00" resultid="7984" heatid="10739" lane="3" entrytime="00:01:10.24" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Guilherme Ballatka" birthdate="2007-06-24" gender="M" nation="BRA" license="398616" swrid="5697228" athleteid="8378" externalid="398616">
              <RESULTS>
                <RESULT eventid="1071" points="438" swimtime="00:02:27.29" resultid="8379" heatid="10478" lane="5" entrytime="00:02:27.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                    <SPLIT distance="100" swimtime="00:01:11.31" />
                    <SPLIT distance="150" swimtime="00:01:49.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="494" swimtime="00:00:58.67" resultid="8380" heatid="10548" lane="7" entrytime="00:01:00.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="516" swimtime="00:00:26.06" resultid="8381" heatid="10626" lane="0" entrytime="00:00:26.04" entrycourse="LCM" />
                <RESULT eventid="1305" points="493" swimtime="00:00:29.80" resultid="8382" heatid="10687" lane="9" entrytime="00:00:30.33" entrycourse="LCM" />
                <RESULT eventid="1373" points="482" swimtime="00:01:05.77" resultid="8383" heatid="10741" lane="7" entrytime="00:01:05.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Wolf Macedo" birthdate="2012-01-27" gender="F" nation="BRA" license="369277" swrid="5602592" athleteid="8202" externalid="369277">
              <RESULTS>
                <RESULT eventid="1079" points="285" swimtime="00:03:28.91" resultid="8203" heatid="10481" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.42" />
                    <SPLIT distance="100" swimtime="00:01:42.62" />
                    <SPLIT distance="150" swimtime="00:02:37.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="441" swimtime="00:01:07.92" resultid="8204" heatid="10532" lane="8" entrytime="00:01:06.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="360" swimtime="00:06:11.62" resultid="8205" heatid="10519" lane="9" entrytime="00:06:24.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                    <SPLIT distance="100" swimtime="00:01:26.46" />
                    <SPLIT distance="150" swimtime="00:02:14.71" />
                    <SPLIT distance="200" swimtime="00:03:03.14" />
                    <SPLIT distance="250" swimtime="00:03:58.48" />
                    <SPLIT distance="300" swimtime="00:04:53.44" />
                    <SPLIT distance="350" swimtime="00:05:33.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="430" swimtime="00:00:31.27" resultid="8206" heatid="10604" lane="8" entrytime="00:00:32.34" entrycourse="LCM" />
                <RESULT eventid="1281" points="456" swimtime="00:02:25.76" resultid="8207" heatid="10657" lane="1" entrytime="00:02:29.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                    <SPLIT distance="100" swimtime="00:01:10.83" />
                    <SPLIT distance="150" swimtime="00:01:49.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="330" swimtime="00:01:19.82" resultid="8208" heatid="10701" lane="0" entrytime="00:01:23.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Artigas Pinheiro" birthdate="2011-08-25" gender="M" nation="BRA" license="377040" swrid="5588535" athleteid="8277" externalid="377040">
              <RESULTS>
                <RESULT eventid="1123" points="385" swimtime="00:10:20.96" resultid="8278" heatid="10516" lane="3" entrytime="00:10:56.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                    <SPLIT distance="100" swimtime="00:01:14.25" />
                    <SPLIT distance="150" swimtime="00:01:52.96" />
                    <SPLIT distance="200" swimtime="00:02:32.49" />
                    <SPLIT distance="250" swimtime="00:03:12.19" />
                    <SPLIT distance="300" swimtime="00:03:51.67" />
                    <SPLIT distance="350" swimtime="00:04:31.66" />
                    <SPLIT distance="400" swimtime="00:05:11.34" />
                    <SPLIT distance="450" swimtime="00:05:51.09" />
                    <SPLIT distance="500" swimtime="00:06:30.69" />
                    <SPLIT distance="550" swimtime="00:07:09.60" />
                    <SPLIT distance="600" swimtime="00:07:48.81" />
                    <SPLIT distance="650" swimtime="00:08:27.78" />
                    <SPLIT distance="700" swimtime="00:09:06.49" />
                    <SPLIT distance="750" swimtime="00:09:44.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="408" swimtime="00:02:49.05" resultid="8279" heatid="10491" lane="7" entrytime="00:02:48.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.73" />
                    <SPLIT distance="100" swimtime="00:01:23.10" />
                    <SPLIT distance="150" swimtime="00:02:07.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="394" swimtime="00:19:47.27" resultid="8280" heatid="10638" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                    <SPLIT distance="100" swimtime="00:01:13.53" />
                    <SPLIT distance="150" swimtime="00:01:52.75" />
                    <SPLIT distance="200" swimtime="00:02:32.49" />
                    <SPLIT distance="250" swimtime="00:03:12.60" />
                    <SPLIT distance="300" swimtime="00:03:52.35" />
                    <SPLIT distance="350" swimtime="00:04:31.82" />
                    <SPLIT distance="400" swimtime="00:05:12.06" />
                    <SPLIT distance="450" swimtime="00:05:51.72" />
                    <SPLIT distance="500" swimtime="00:06:31.53" />
                    <SPLIT distance="550" swimtime="00:07:11.08" />
                    <SPLIT distance="600" swimtime="00:07:51.38" />
                    <SPLIT distance="650" swimtime="00:08:31.07" />
                    <SPLIT distance="700" swimtime="00:09:11.27" />
                    <SPLIT distance="750" swimtime="00:09:51.24" />
                    <SPLIT distance="800" swimtime="00:10:31.40" />
                    <SPLIT distance="850" swimtime="00:11:10.84" />
                    <SPLIT distance="900" swimtime="00:11:51.12" />
                    <SPLIT distance="950" swimtime="00:12:31.03" />
                    <SPLIT distance="1000" swimtime="00:13:11.38" />
                    <SPLIT distance="1050" swimtime="00:13:51.08" />
                    <SPLIT distance="1100" swimtime="00:14:31.38" />
                    <SPLIT distance="1150" swimtime="00:15:11.11" />
                    <SPLIT distance="1200" swimtime="00:15:51.39" />
                    <SPLIT distance="1250" swimtime="00:16:30.71" />
                    <SPLIT distance="1300" swimtime="00:17:11.21" />
                    <SPLIT distance="1350" swimtime="00:17:51.19" />
                    <SPLIT distance="1400" swimtime="00:18:31.24" />
                    <SPLIT distance="1450" swimtime="00:19:09.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="344" swimtime="00:01:21.13" resultid="8281" heatid="10595" lane="5" entrytime="00:01:21.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="353" swimtime="00:02:41.30" resultid="8282" heatid="10648" lane="1" entrytime="00:02:51.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.31" />
                    <SPLIT distance="100" swimtime="00:01:20.59" />
                    <SPLIT distance="150" swimtime="00:02:04.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="393" swimtime="00:05:00.42" resultid="8283" heatid="10719" lane="2" entrytime="00:05:27.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                    <SPLIT distance="100" swimtime="00:01:10.75" />
                    <SPLIT distance="150" swimtime="00:01:48.77" />
                    <SPLIT distance="200" swimtime="00:02:27.67" />
                    <SPLIT distance="250" swimtime="00:03:06.50" />
                    <SPLIT distance="300" swimtime="00:03:45.34" />
                    <SPLIT distance="350" swimtime="00:04:23.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="David Cella" birthdate="2008-02-17" gender="M" nation="BRA" license="341107" swrid="5634581" athleteid="8337" externalid="341107">
              <RESULTS>
                <RESULT eventid="1187" points="577" swimtime="00:00:31.16" resultid="8338" heatid="10575" lane="6" entrytime="00:00:30.11" entrycourse="LCM" />
                <RESULT eventid="1155" points="644" swimtime="00:00:53.73" resultid="8339" heatid="10552" lane="6" entrytime="00:00:52.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="594" swimtime="00:00:24.87" resultid="8340" heatid="10628" lane="6" entrytime="00:00:24.11" entrycourse="LCM" />
                <RESULT eventid="1219" status="WDR" swimtime="00:00:00.00" resultid="8341" heatid="10598" lane="6" entrytime="00:01:11.80" entrycourse="LCM" />
                <RESULT eventid="1289" points="494" swimtime="00:02:09.02" resultid="8342" heatid="10664" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.48" />
                    <SPLIT distance="100" swimtime="00:01:00.33" />
                    <SPLIT distance="150" swimtime="00:01:35.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="532" swimtime="00:01:03.68" resultid="8343" heatid="10742" lane="1" entrytime="00:01:03.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Karam Barbosa Lima" birthdate="2012-12-11" gender="F" nation="BRA" license="376956" swrid="5588758" athleteid="8254" externalid="376956">
              <RESULTS>
                <RESULT eventid="1063" points="340" swimtime="00:02:56.38" resultid="8255" heatid="10471" lane="2" entrytime="00:02:53.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.87" />
                    <SPLIT distance="100" swimtime="00:01:25.82" />
                    <SPLIT distance="150" swimtime="00:02:11.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="366" swimtime="00:01:12.28" resultid="8256" heatid="10528" lane="2" entrytime="00:01:12.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 9:40)" eventid="1227" status="DSQ" swimtime="00:00:32.55" resultid="8257" heatid="10604" lane="6" entrytime="00:00:32.09" entrycourse="LCM" />
                <RESULT eventid="1281" points="351" swimtime="00:02:39.09" resultid="8258" heatid="10653" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                    <SPLIT distance="100" swimtime="00:01:14.92" />
                    <SPLIT distance="150" swimtime="00:01:57.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="356" swimtime="00:01:20.55" resultid="8259" heatid="10730" lane="0" entrytime="00:01:20.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joshua" lastname="Gomide Capraro" birthdate="2009-01-18" gender="M" nation="BRA" license="339030" swrid="5600177" athleteid="7846" externalid="339030">
              <RESULTS>
                <RESULT eventid="1103" status="DNS" swimtime="00:00:00.00" resultid="7847" heatid="10507" lane="7" entrytime="00:00:28.59" entrycourse="LCM" />
                <RESULT eventid="1155" status="DNS" swimtime="00:00:00.00" resultid="7848" heatid="10552" lane="0" entrytime="00:00:54.26" entrycourse="LCM" />
                <RESULT eventid="1235" status="DNS" swimtime="00:00:00.00" resultid="7849" heatid="10628" lane="0" entrytime="00:00:24.57" entrycourse="LCM" />
                <RESULT eventid="1289" status="DNS" swimtime="00:00:00.00" resultid="7850" heatid="10673" lane="4" entrytime="00:02:02.43" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Lazzarotti Matias" birthdate="2012-03-19" gender="F" nation="BRA" license="391026" swrid="5602552" athleteid="8314" externalid="391026">
              <RESULTS>
                <RESULT eventid="1063" points="384" swimtime="00:02:49.34" resultid="8315" heatid="10471" lane="3" entrytime="00:02:52.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                    <SPLIT distance="100" swimtime="00:01:23.77" />
                    <SPLIT distance="150" swimtime="00:02:07.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="401" swimtime="00:01:10.08" resultid="8316" heatid="10529" lane="6" entrytime="00:01:10.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="286" swimtime="00:01:37.33" resultid="8317" heatid="10584" lane="4" entrytime="00:01:36.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="418" swimtime="00:02:30.00" resultid="8318" heatid="10656" lane="5" entrytime="00:02:31.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                    <SPLIT distance="100" swimtime="00:01:13.91" />
                    <SPLIT distance="150" swimtime="00:01:53.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="364" swimtime="00:05:29.46" resultid="8319" heatid="10714" lane="6" entrytime="00:05:16.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="100" swimtime="00:01:16.43" />
                    <SPLIT distance="150" swimtime="00:01:59.03" />
                    <SPLIT distance="200" swimtime="00:02:41.22" />
                    <SPLIT distance="250" swimtime="00:03:23.64" />
                    <SPLIT distance="300" swimtime="00:04:06.28" />
                    <SPLIT distance="350" swimtime="00:04:48.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="389" swimtime="00:01:18.22" resultid="8320" heatid="10730" lane="2" entrytime="00:01:18.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Galvao" birthdate="2011-03-11" gender="M" nation="BRA" license="381989" swrid="5602541" athleteid="8292" externalid="381989">
              <RESULTS>
                <RESULT eventid="1103" points="228" swimtime="00:00:36.44" resultid="8293" heatid="10500" lane="9" />
                <RESULT eventid="1171" points="178" swimtime="00:03:15.93" resultid="8294" heatid="10555" lane="4" entrytime="00:03:21.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.81" />
                    <SPLIT distance="100" swimtime="00:01:34.26" />
                    <SPLIT distance="150" swimtime="00:02:28.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="344" swimtime="00:01:06.16" resultid="8295" heatid="10544" lane="6" entrytime="00:01:06.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="318" swimtime="00:00:30.63" resultid="8296" heatid="10617" lane="5" entrytime="00:00:31.01" entrycourse="LCM" />
                <RESULT eventid="1341" points="206" swimtime="00:01:23.65" resultid="8297" heatid="10705" lane="5" entrytime="00:01:25.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Cabrera Cirino" birthdate="2011-01-28" gender="M" nation="BRA" license="369531" swrid="5588569" athleteid="8235" externalid="369531">
              <RESULTS>
                <RESULT eventid="1123" points="471" swimtime="00:09:40.99" resultid="8236" heatid="10514" lane="2" entrytime="00:09:46.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                    <SPLIT distance="100" swimtime="00:01:08.41" />
                    <SPLIT distance="150" swimtime="00:01:44.20" />
                    <SPLIT distance="200" swimtime="00:02:20.18" />
                    <SPLIT distance="250" swimtime="00:02:56.85" />
                    <SPLIT distance="300" swimtime="00:03:33.73" />
                    <SPLIT distance="350" swimtime="00:04:10.78" />
                    <SPLIT distance="400" swimtime="00:04:47.26" />
                    <SPLIT distance="450" swimtime="00:05:24.17" />
                    <SPLIT distance="500" swimtime="00:06:00.64" />
                    <SPLIT distance="550" swimtime="00:06:37.66" />
                    <SPLIT distance="600" swimtime="00:07:14.81" />
                    <SPLIT distance="650" swimtime="00:07:52.28" />
                    <SPLIT distance="700" swimtime="00:08:28.90" />
                    <SPLIT distance="750" swimtime="00:09:05.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="427" swimtime="00:02:28.52" resultid="8237" heatid="10479" lane="1" entrytime="00:02:26.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                    <SPLIT distance="100" swimtime="00:01:11.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="490" swimtime="00:00:58.82" resultid="8238" heatid="10549" lane="7" entrytime="00:00:58.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="506" swimtime="00:00:26.24" resultid="8239" heatid="10624" lane="5" entrytime="00:00:26.96" entrycourse="LCM" />
                <RESULT eventid="1289" points="515" swimtime="00:02:07.25" resultid="8240" heatid="10672" lane="8" entrytime="00:02:09.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.16" />
                    <SPLIT distance="100" swimtime="00:01:01.86" />
                    <SPLIT distance="150" swimtime="00:01:35.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="506" swimtime="00:04:36.11" resultid="8241" heatid="10723" lane="1" entrytime="00:04:36.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.36" />
                    <SPLIT distance="100" swimtime="00:01:04.13" />
                    <SPLIT distance="150" swimtime="00:01:38.30" />
                    <SPLIT distance="200" swimtime="00:02:13.77" />
                    <SPLIT distance="250" swimtime="00:02:49.21" />
                    <SPLIT distance="300" swimtime="00:03:25.24" />
                    <SPLIT distance="350" swimtime="00:04:01.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luana" lastname="Zeclhynski Silva" birthdate="2006-09-14" gender="F" nation="BRA" license="330727" swrid="5600283" athleteid="7832" externalid="330727" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1297" points="680" swimtime="00:00:30.53" resultid="7833" heatid="10680" lane="4" entrytime="00:00:30.32" entrycourse="LCM" />
                <RESULT eventid="1365" points="656" swimtime="00:01:05.75" resultid="7834" heatid="10732" lane="4" entrytime="00:01:05.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Presiazniuk" birthdate="2010-10-14" gender="M" nation="BRA" license="356353" swrid="5600237" athleteid="7999" externalid="356353">
              <RESULTS>
                <RESULT eventid="1071" points="449" swimtime="00:02:26.14" resultid="8000" heatid="10478" lane="4" entrytime="00:02:27.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                    <SPLIT distance="100" swimtime="00:01:11.58" />
                    <SPLIT distance="150" swimtime="00:01:49.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="509" swimtime="00:00:58.11" resultid="8001" heatid="10549" lane="3" entrytime="00:00:58.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="469" swimtime="00:00:26.90" resultid="8002" heatid="10623" lane="3" entrytime="00:00:27.51" entrycourse="LCM" />
                <RESULT eventid="1273" points="394" swimtime="00:02:35.44" resultid="8003" heatid="10649" lane="6" entrytime="00:02:40.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                    <SPLIT distance="100" swimtime="00:01:12.23" />
                    <SPLIT distance="150" swimtime="00:02:03.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="492" swimtime="00:02:09.19" resultid="8004" heatid="10672" lane="9" entrytime="00:02:09.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.67" />
                    <SPLIT distance="100" swimtime="00:01:02.82" />
                    <SPLIT distance="150" swimtime="00:01:36.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="445" swimtime="00:01:07.58" resultid="8005" heatid="10740" lane="7" entrytime="00:01:08.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Iglesias Vargas" birthdate="2009-01-11" gender="M" nation="BRA" license="324792" swrid="5600189" athleteid="7884" externalid="324792">
              <RESULTS>
                <RESULT eventid="1123" points="536" swimtime="00:09:16.45" resultid="7885" heatid="10513" lane="1" entrytime="00:09:11.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.26" />
                    <SPLIT distance="100" swimtime="00:01:05.15" />
                    <SPLIT distance="150" swimtime="00:01:39.42" />
                    <SPLIT distance="200" swimtime="00:02:13.83" />
                    <SPLIT distance="250" swimtime="00:02:48.41" />
                    <SPLIT distance="300" swimtime="00:03:23.18" />
                    <SPLIT distance="350" swimtime="00:03:57.92" />
                    <SPLIT distance="400" swimtime="00:04:32.98" />
                    <SPLIT distance="450" swimtime="00:05:07.98" />
                    <SPLIT distance="500" swimtime="00:05:43.54" />
                    <SPLIT distance="550" swimtime="00:06:19.09" />
                    <SPLIT distance="600" swimtime="00:06:54.91" />
                    <SPLIT distance="650" swimtime="00:07:30.88" />
                    <SPLIT distance="700" swimtime="00:08:06.60" />
                    <SPLIT distance="750" swimtime="00:08:42.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="577" swimtime="00:00:55.72" resultid="7886" heatid="10551" lane="8" entrytime="00:00:56.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="607" swimtime="00:02:00.44" resultid="7887" heatid="10674" lane="9" entrytime="00:02:01.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.26" />
                    <SPLIT distance="100" swimtime="00:00:57.14" />
                    <SPLIT distance="150" swimtime="00:01:28.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="588" swimtime="00:04:22.66" resultid="7888" heatid="10724" lane="7" entrytime="00:04:23.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.65" />
                    <SPLIT distance="100" swimtime="00:01:01.89" />
                    <SPLIT distance="150" swimtime="00:01:34.96" />
                    <SPLIT distance="200" swimtime="00:02:08.73" />
                    <SPLIT distance="250" swimtime="00:02:42.92" />
                    <SPLIT distance="300" swimtime="00:03:16.93" />
                    <SPLIT distance="350" swimtime="00:03:50.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Petraglia" birthdate="2012-03-28" gender="M" nation="BRA" license="369282" swrid="5602569" athleteid="8228" externalid="369282">
              <RESULTS>
                <RESULT eventid="1071" points="263" swimtime="00:02:54.62" resultid="8229" heatid="10476" lane="9" entrytime="00:02:59.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.14" />
                    <SPLIT distance="100" swimtime="00:01:25.17" />
                    <SPLIT distance="150" swimtime="00:02:10.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="208" swimtime="00:00:43.77" resultid="8230" heatid="10571" lane="7" entrytime="00:00:43.53" entrycourse="LCM" />
                <RESULT eventid="1155" points="257" swimtime="00:01:12.96" resultid="8231" heatid="10535" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="192" swimtime="00:01:38.46" resultid="8232" heatid="10592" lane="3" entrytime="00:01:39.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" status="DNS" swimtime="00:00:00.00" resultid="8233" heatid="10663" lane="2" />
                <RESULT eventid="1373" points="233" swimtime="00:01:23.83" resultid="8234" heatid="10736" lane="8" entrytime="00:01:25.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Rocha" birthdate="2011-08-25" gender="F" nation="BRA" license="366904" swrid="5602578" athleteid="8083" externalid="366904">
              <RESULTS>
                <RESULT eventid="1063" points="388" swimtime="00:02:48.72" resultid="8084" heatid="10472" lane="0" entrytime="00:02:48.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                    <SPLIT distance="100" swimtime="00:01:23.47" />
                    <SPLIT distance="150" swimtime="00:02:06.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="477" swimtime="00:01:06.16" resultid="8085" heatid="10533" lane="8" entrytime="00:01:05.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="457" swimtime="00:00:30.65" resultid="8086" heatid="10607" lane="7" entrytime="00:00:30.29" entrycourse="LCM" />
                <RESULT eventid="1281" points="425" swimtime="00:02:29.27" resultid="8087" heatid="10659" lane="8" entrytime="00:02:23.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.88" />
                    <SPLIT distance="100" swimtime="00:01:10.54" />
                    <SPLIT distance="150" swimtime="00:01:50.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="414" swimtime="00:05:15.58" resultid="8088" heatid="10715" lane="6" entrytime="00:05:06.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                    <SPLIT distance="100" swimtime="00:01:13.69" />
                    <SPLIT distance="150" swimtime="00:01:53.40" />
                    <SPLIT distance="200" swimtime="00:02:33.79" />
                    <SPLIT distance="250" swimtime="00:03:14.27" />
                    <SPLIT distance="300" swimtime="00:03:55.06" />
                    <SPLIT distance="350" swimtime="00:04:35.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="358" swimtime="00:01:20.39" resultid="8089" heatid="10730" lane="3" entrytime="00:01:18.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Zaroni" birthdate="2010-03-03" gender="F" nation="BRA" license="356345" swrid="5600282" athleteid="7871" externalid="356345">
              <RESULTS>
                <RESULT eventid="1095" points="351" swimtime="00:00:34.63" resultid="7872" heatid="10497" lane="9" entrytime="00:00:36.35" entrycourse="LCM" />
                <RESULT eventid="1079" points="503" swimtime="00:02:52.92" resultid="7873" heatid="10486" lane="6" entrytime="00:02:53.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.51" />
                    <SPLIT distance="100" swimtime="00:01:24.89" />
                    <SPLIT distance="150" swimtime="00:02:09.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="503" swimtime="00:01:05.01" resultid="7874" heatid="10532" lane="3" entrytime="00:01:05.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="462" swimtime="00:01:22.92" resultid="7875" heatid="10588" lane="2" entrytime="00:01:22.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="379" swimtime="00:00:37.09" resultid="7876" heatid="10676" lane="2" />
                <RESULT eventid="1265" points="469" swimtime="00:02:42.32" resultid="7877" heatid="10643" lane="7" entrytime="00:02:45.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                    <SPLIT distance="100" swimtime="00:01:18.88" />
                    <SPLIT distance="150" swimtime="00:02:04.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Salomao" birthdate="2012-05-07" gender="M" nation="BRA" license="369261" swrid="5602581" athleteid="8135" externalid="369261">
              <RESULTS>
                <RESULT eventid="1123" points="296" swimtime="00:11:18.03" resultid="8136" heatid="10517" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                    <SPLIT distance="100" swimtime="00:01:17.85" />
                    <SPLIT distance="150" swimtime="00:01:59.56" />
                    <SPLIT distance="200" swimtime="00:02:43.07" />
                    <SPLIT distance="250" swimtime="00:03:25.57" />
                    <SPLIT distance="300" swimtime="00:04:07.95" />
                    <SPLIT distance="350" swimtime="00:04:50.32" />
                    <SPLIT distance="400" swimtime="00:05:33.59" />
                    <SPLIT distance="450" swimtime="00:06:17.28" />
                    <SPLIT distance="500" swimtime="00:06:59.88" />
                    <SPLIT distance="550" swimtime="00:07:42.05" />
                    <SPLIT distance="600" swimtime="00:08:26.21" />
                    <SPLIT distance="650" swimtime="00:09:10.52" />
                    <SPLIT distance="700" swimtime="00:09:53.50" />
                    <SPLIT distance="750" swimtime="00:10:37.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="245" swimtime="00:02:58.64" resultid="8137" heatid="10475" lane="4" entrytime="00:03:09.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.18" />
                    <SPLIT distance="100" swimtime="00:01:27.03" />
                    <SPLIT distance="150" swimtime="00:02:14.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="281" swimtime="00:00:31.92" resultid="8138" heatid="10615" lane="2" entrytime="00:00:32.53" entrycourse="LCM" />
                <RESULT eventid="1289" points="296" swimtime="00:02:33.05" resultid="8139" heatid="10666" lane="6" entrytime="00:02:35.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.03" />
                    <SPLIT distance="100" swimtime="00:01:13.75" />
                    <SPLIT distance="150" swimtime="00:01:53.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="316" swimtime="00:05:22.88" resultid="8140" heatid="10719" lane="7" entrytime="00:05:28.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                    <SPLIT distance="100" swimtime="00:01:16.34" />
                    <SPLIT distance="150" swimtime="00:01:57.49" />
                    <SPLIT distance="200" swimtime="00:02:39.88" />
                    <SPLIT distance="250" swimtime="00:03:21.06" />
                    <SPLIT distance="300" swimtime="00:04:03.43" />
                    <SPLIT distance="350" swimtime="00:04:43.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="181" swimtime="00:01:31.13" resultid="8141" heatid="10734" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Antunes Saboia" birthdate="2012-06-28" gender="M" nation="BRA" license="369278" swrid="5602511" athleteid="8209" externalid="369278">
              <RESULTS>
                <RESULT eventid="1087" points="314" swimtime="00:03:04.54" resultid="8210" heatid="10489" lane="3" entrytime="00:03:04.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.59" />
                    <SPLIT distance="100" swimtime="00:01:29.14" />
                    <SPLIT distance="150" swimtime="00:02:17.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="323" swimtime="00:01:07.61" resultid="8211" heatid="10542" lane="1" entrytime="00:01:09.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="306" swimtime="00:01:24.32" resultid="8212" heatid="10595" lane="9" entrytime="00:01:25.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 6.5 - Não terminou a prova enquanto estava de costas.&#10;&#10;&#10;&#10;&#10;&#10;&#10;  (Horário: 16:43), Na volta dos 100m (Costas, Medley Individual)." eventid="1273" status="DSQ" swimtime="00:02:51.88" resultid="8213" heatid="10648" lane="0" entrytime="00:02:54.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.40" />
                    <SPLIT distance="100" swimtime="00:01:26.33" />
                    <SPLIT distance="150" swimtime="00:02:13.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="214" swimtime="00:01:26.24" resultid="8214" heatid="10736" lane="0" entrytime="00:01:25.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Job Pigatto" birthdate="2012-04-17" gender="M" nation="BRA" license="371100" swrid="5627271" athleteid="8384" externalid="371100">
              <RESULTS>
                <RESULT eventid="1071" points="439" swimtime="00:02:27.16" resultid="8385" heatid="10478" lane="2" entrytime="00:02:30.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                    <SPLIT distance="100" swimtime="00:01:10.10" />
                    <SPLIT distance="150" swimtime="00:01:48.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="471" swimtime="00:00:59.60" resultid="8386" heatid="10546" lane="0" entrytime="00:01:03.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="448" swimtime="00:00:27.31" resultid="8387" heatid="10622" lane="7" entrytime="00:00:28.09" entrycourse="LCM" />
                <RESULT eventid="1289" points="462" swimtime="00:02:11.93" resultid="8388" heatid="10671" lane="0" entrytime="00:02:15.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.23" />
                    <SPLIT distance="100" swimtime="00:01:02.33" />
                    <SPLIT distance="150" swimtime="00:01:37.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="416" swimtime="00:01:09.09" resultid="8389" heatid="10739" lane="4" entrytime="00:01:09.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Viera Correa" birthdate="2012-03-07" gender="M" nation="BRA" license="369269" swrid="5602590" athleteid="8162" externalid="369269">
              <RESULTS>
                <RESULT eventid="1123" points="346" swimtime="00:10:43.75" resultid="8163" heatid="10517" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.08" />
                    <SPLIT distance="100" swimtime="00:01:16.01" />
                    <SPLIT distance="150" swimtime="00:01:56.51" />
                    <SPLIT distance="200" swimtime="00:02:37.63" />
                    <SPLIT distance="250" swimtime="00:03:17.85" />
                    <SPLIT distance="300" swimtime="00:03:58.92" />
                    <SPLIT distance="350" swimtime="00:04:39.67" />
                    <SPLIT distance="400" swimtime="00:05:21.07" />
                    <SPLIT distance="450" swimtime="00:06:02.38" />
                    <SPLIT distance="500" swimtime="00:06:43.93" />
                    <SPLIT distance="550" swimtime="00:07:24.47" />
                    <SPLIT distance="600" swimtime="00:08:05.06" />
                    <SPLIT distance="650" swimtime="00:08:46.09" />
                    <SPLIT distance="700" swimtime="00:09:27.15" />
                    <SPLIT distance="750" swimtime="00:10:05.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="295" swimtime="00:02:47.99" resultid="8164" heatid="10476" lane="1" entrytime="00:02:50.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.62" />
                    <SPLIT distance="100" swimtime="00:01:20.36" />
                    <SPLIT distance="150" swimtime="00:02:04.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="363" swimtime="00:01:04.99" resultid="8165" heatid="10544" lane="8" entrytime="00:01:06.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="347" swimtime="00:00:29.73" resultid="8166" heatid="10619" lane="7" entrytime="00:00:29.88" entrycourse="LCM" />
                <RESULT eventid="1289" points="354" swimtime="00:02:24.13" resultid="8167" heatid="10667" lane="3" entrytime="00:02:28.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                    <SPLIT distance="100" swimtime="00:01:08.35" />
                    <SPLIT distance="150" swimtime="00:01:46.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="278" swimtime="00:01:19.05" resultid="8168" heatid="10736" lane="6" entrytime="00:01:21.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcelo" lastname="Vanhazebrouck" birthdate="2010-01-09" gender="M" nation="BRA" license="339043" swrid="5600269" athleteid="7971" externalid="339043">
              <RESULTS>
                <RESULT eventid="1103" points="343" swimtime="00:00:31.79" resultid="7972" heatid="10505" lane="6" entrytime="00:00:31.37" entrycourse="LCM" />
                <RESULT eventid="1187" points="360" swimtime="00:00:36.46" resultid="7973" heatid="10569" lane="5" />
                <RESULT eventid="1155" points="429" swimtime="00:01:01.51" resultid="7974" heatid="10548" lane="2" entrytime="00:01:00.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="420" swimtime="00:00:27.92" resultid="7975" heatid="10623" lane="6" entrytime="00:00:27.57" entrycourse="LCM" />
                <RESULT eventid="1219" points="325" swimtime="00:01:22.67" resultid="7976" heatid="10595" lane="1" entrytime="00:01:23.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="399" swimtime="00:02:18.46" resultid="7977" heatid="10671" lane="9" entrytime="00:02:15.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.87" />
                    <SPLIT distance="100" swimtime="00:01:05.73" />
                    <SPLIT distance="150" swimtime="00:01:41.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabrizio" lastname="Bulla Lanaro" birthdate="2009-08-28" gender="M" nation="BRA" license="344303" swrid="5559846" athleteid="8373" externalid="344303">
              <RESULTS>
                <RESULT eventid="1103" points="498" swimtime="00:00:28.08" resultid="8374" heatid="10508" lane="0" entrytime="00:00:27.60" entrycourse="LCM" />
                <RESULT eventid="1187" points="556" swimtime="00:00:31.54" resultid="8375" heatid="10569" lane="2" />
                <RESULT eventid="1219" points="533" swimtime="00:01:10.13" resultid="8376" heatid="10598" lane="5" entrytime="00:01:09.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="501" swimtime="00:01:02.23" resultid="8377" heatid="10710" lane="3" entrytime="00:01:01.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Kraemer Geremia" birthdate="2011-07-20" gender="F" nation="BRA" license="366908" swrid="5588763" athleteid="8104" externalid="366908">
              <RESULTS>
                <RESULT eventid="1115" points="404" swimtime="00:20:44.53" resultid="8105" heatid="10511" lane="7" entrytime="00:20:00.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                    <SPLIT distance="100" swimtime="00:01:15.62" />
                    <SPLIT distance="150" swimtime="00:01:55.91" />
                    <SPLIT distance="200" swimtime="00:02:36.96" />
                    <SPLIT distance="250" swimtime="00:03:18.17" />
                    <SPLIT distance="300" swimtime="00:04:00.14" />
                    <SPLIT distance="350" swimtime="00:04:41.23" />
                    <SPLIT distance="400" swimtime="00:05:23.27" />
                    <SPLIT distance="450" swimtime="00:06:04.68" />
                    <SPLIT distance="500" swimtime="00:06:46.85" />
                    <SPLIT distance="550" swimtime="00:07:29.09" />
                    <SPLIT distance="600" swimtime="00:08:11.37" />
                    <SPLIT distance="650" swimtime="00:08:53.66" />
                    <SPLIT distance="700" swimtime="00:09:36.96" />
                    <SPLIT distance="750" swimtime="00:10:20.26" />
                    <SPLIT distance="800" swimtime="00:11:03.01" />
                    <SPLIT distance="850" swimtime="00:11:46.49" />
                    <SPLIT distance="900" swimtime="00:12:29.10" />
                    <SPLIT distance="950" swimtime="00:13:11.63" />
                    <SPLIT distance="1000" swimtime="00:13:53.76" />
                    <SPLIT distance="1050" swimtime="00:14:35.71" />
                    <SPLIT distance="1100" swimtime="00:15:17.77" />
                    <SPLIT distance="1150" swimtime="00:15:59.93" />
                    <SPLIT distance="1200" swimtime="00:16:41.63" />
                    <SPLIT distance="1250" swimtime="00:17:23.16" />
                    <SPLIT distance="1300" swimtime="00:18:03.87" />
                    <SPLIT distance="1350" swimtime="00:18:44.66" />
                    <SPLIT distance="1400" swimtime="00:19:25.20" />
                    <SPLIT distance="1450" swimtime="00:20:05.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="442" swimtime="00:02:41.62" resultid="8106" heatid="10473" lane="1" entrytime="00:02:38.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                    <SPLIT distance="100" swimtime="00:01:18.68" />
                    <SPLIT distance="150" swimtime="00:01:59.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="485" swimtime="00:01:05.79" resultid="8107" heatid="10533" lane="7" entrytime="00:01:05.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="456" swimtime="00:10:29.81" resultid="8108" heatid="10632" lane="5" entrytime="00:10:14.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                    <SPLIT distance="100" swimtime="00:01:11.52" />
                    <SPLIT distance="150" swimtime="00:01:50.62" />
                    <SPLIT distance="200" swimtime="00:02:30.14" />
                    <SPLIT distance="250" swimtime="00:03:09.75" />
                    <SPLIT distance="300" swimtime="00:03:49.67" />
                    <SPLIT distance="350" swimtime="00:04:29.44" />
                    <SPLIT distance="400" swimtime="00:05:08.97" />
                    <SPLIT distance="450" swimtime="00:05:48.99" />
                    <SPLIT distance="500" swimtime="00:06:28.83" />
                    <SPLIT distance="550" swimtime="00:07:09.20" />
                    <SPLIT distance="600" swimtime="00:07:49.63" />
                    <SPLIT distance="650" swimtime="00:08:30.06" />
                    <SPLIT distance="700" swimtime="00:09:10.65" />
                    <SPLIT distance="750" swimtime="00:09:50.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="478" swimtime="00:02:23.51" resultid="8109" heatid="10659" lane="6" entrytime="00:02:22.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                    <SPLIT distance="100" swimtime="00:01:09.89" />
                    <SPLIT distance="150" swimtime="00:01:47.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="444" swimtime="00:05:08.48" resultid="8110" heatid="10716" lane="2" entrytime="00:04:58.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                    <SPLIT distance="100" swimtime="00:01:12.30" />
                    <SPLIT distance="150" swimtime="00:01:51.41" />
                    <SPLIT distance="200" swimtime="00:02:31.29" />
                    <SPLIT distance="250" swimtime="00:03:10.94" />
                    <SPLIT distance="300" swimtime="00:03:50.89" />
                    <SPLIT distance="350" swimtime="00:04:29.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Almeida Pinheiro" birthdate="2005-06-29" gender="M" nation="BRA" license="331635" swrid="5330117" athleteid="8406" externalid="331635">
              <RESULTS>
                <RESULT eventid="1171" points="678" swimtime="00:02:05.60" resultid="8407" heatid="10558" lane="4" entrytime="00:02:03.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                    <SPLIT distance="100" swimtime="00:00:59.04" />
                    <SPLIT distance="150" swimtime="00:01:31.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="672" swimtime="00:01:56.40" resultid="8408" heatid="10674" lane="3" entrytime="00:01:56.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.77" />
                    <SPLIT distance="100" swimtime="00:00:56.44" />
                    <SPLIT distance="150" swimtime="00:01:26.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Mattioli" birthdate="2011-10-22" gender="F" nation="BRA" license="366896" swrid="5602559" athleteid="8062" externalid="366896">
              <RESULTS>
                <RESULT eventid="1115" points="431" swimtime="00:20:18.04" resultid="8063" heatid="10511" lane="2" entrytime="00:19:57.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.46" />
                    <SPLIT distance="100" swimtime="00:01:15.62" />
                    <SPLIT distance="150" swimtime="00:01:56.58" />
                    <SPLIT distance="200" swimtime="00:02:38.47" />
                    <SPLIT distance="250" swimtime="00:03:19.17" />
                    <SPLIT distance="300" swimtime="00:04:00.24" />
                    <SPLIT distance="350" swimtime="00:04:41.51" />
                    <SPLIT distance="400" swimtime="00:05:23.19" />
                    <SPLIT distance="450" swimtime="00:06:04.03" />
                    <SPLIT distance="500" swimtime="00:06:44.83" />
                    <SPLIT distance="550" swimtime="00:07:25.49" />
                    <SPLIT distance="600" swimtime="00:08:06.74" />
                    <SPLIT distance="650" swimtime="00:08:47.85" />
                    <SPLIT distance="700" swimtime="00:09:28.35" />
                    <SPLIT distance="750" swimtime="00:10:09.96" />
                    <SPLIT distance="800" swimtime="00:10:51.20" />
                    <SPLIT distance="850" swimtime="00:11:31.82" />
                    <SPLIT distance="900" swimtime="00:12:13.44" />
                    <SPLIT distance="950" swimtime="00:12:55.54" />
                    <SPLIT distance="1000" swimtime="00:13:37.21" />
                    <SPLIT distance="1050" swimtime="00:14:18.07" />
                    <SPLIT distance="1100" swimtime="00:14:58.76" />
                    <SPLIT distance="1150" swimtime="00:15:39.52" />
                    <SPLIT distance="1200" swimtime="00:16:20.46" />
                    <SPLIT distance="1250" swimtime="00:17:00.85" />
                    <SPLIT distance="1300" swimtime="00:17:41.85" />
                    <SPLIT distance="1350" swimtime="00:18:22.20" />
                    <SPLIT distance="1400" swimtime="00:19:02.43" />
                    <SPLIT distance="1450" swimtime="00:19:41.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="520" swimtime="00:02:51.02" resultid="8064" heatid="10486" lane="3" entrytime="00:02:51.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.87" />
                    <SPLIT distance="100" swimtime="00:01:22.71" />
                    <SPLIT distance="150" swimtime="00:02:07.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="451" swimtime="00:05:44.73" resultid="8065" heatid="10518" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.12" />
                    <SPLIT distance="100" swimtime="00:01:26.20" />
                    <SPLIT distance="150" swimtime="00:02:12.82" />
                    <SPLIT distance="200" swimtime="00:02:59.96" />
                    <SPLIT distance="250" swimtime="00:03:44.91" />
                    <SPLIT distance="300" swimtime="00:04:30.21" />
                    <SPLIT distance="350" swimtime="00:05:08.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="483" swimtime="00:10:17.51" resultid="8066" heatid="10632" lane="7" entrytime="00:10:34.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                    <SPLIT distance="100" swimtime="00:01:12.43" />
                    <SPLIT distance="150" swimtime="00:01:52.07" />
                    <SPLIT distance="200" swimtime="00:02:31.50" />
                    <SPLIT distance="250" swimtime="00:03:10.86" />
                    <SPLIT distance="300" swimtime="00:03:50.56" />
                    <SPLIT distance="350" swimtime="00:04:29.75" />
                    <SPLIT distance="400" swimtime="00:05:09.35" />
                    <SPLIT distance="450" swimtime="00:05:47.97" />
                    <SPLIT distance="500" swimtime="00:06:26.74" />
                    <SPLIT distance="550" swimtime="00:07:05.90" />
                    <SPLIT distance="600" swimtime="00:07:45.59" />
                    <SPLIT distance="650" swimtime="00:08:25.00" />
                    <SPLIT distance="700" swimtime="00:09:04.54" />
                    <SPLIT distance="750" swimtime="00:09:42.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="485" swimtime="00:01:21.62" resultid="8067" heatid="10589" lane="0" entrytime="00:01:20.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="473" swimtime="00:02:41.76" resultid="8068" heatid="10643" lane="6" entrytime="00:02:44.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                    <SPLIT distance="100" swimtime="00:01:22.29" />
                    <SPLIT distance="150" swimtime="00:02:07.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Cipriani Presiazniuk" birthdate="2012-07-03" gender="M" nation="BRA" license="369267" swrid="5588594" athleteid="8156" externalid="369267">
              <RESULTS>
                <RESULT eventid="1071" points="268" swimtime="00:02:53.49" resultid="8157" heatid="10476" lane="0" entrytime="00:02:57.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.17" />
                    <SPLIT distance="100" swimtime="00:01:24.89" />
                    <SPLIT distance="150" swimtime="00:02:09.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="306" swimtime="00:01:08.84" resultid="8158" heatid="10541" lane="3" entrytime="00:01:10.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="304" swimtime="00:00:31.07" resultid="8159" heatid="10617" lane="2" entrytime="00:00:31.10" entrycourse="LCM" />
                <RESULT eventid="1289" points="291" swimtime="00:02:33.82" resultid="8160" heatid="10666" lane="9" entrytime="00:02:40.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                    <SPLIT distance="100" swimtime="00:01:14.28" />
                    <SPLIT distance="150" swimtime="00:01:56.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="253" swimtime="00:01:21.50" resultid="8161" heatid="10736" lane="2" entrytime="00:01:21.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cecilia" lastname="Cabrini Vieira" birthdate="2012-02-11" gender="F" nation="BRA" license="376961" swrid="5588571" athleteid="8260" externalid="376961">
              <RESULTS>
                <RESULT eventid="1063" points="418" swimtime="00:02:44.66" resultid="8261" heatid="10471" lane="5" entrytime="00:02:52.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.70" />
                    <SPLIT distance="100" swimtime="00:01:20.47" />
                    <SPLIT distance="150" swimtime="00:02:03.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="521" swimtime="00:01:04.25" resultid="8262" heatid="10532" lane="4" entrytime="00:01:05.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="504" swimtime="00:00:29.65" resultid="8263" heatid="10608" lane="8" entrytime="00:00:29.69" entrycourse="LCM" />
                <RESULT eventid="1281" points="485" swimtime="00:02:22.79" resultid="8264" heatid="10658" lane="0" entrytime="00:02:26.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                    <SPLIT distance="100" swimtime="00:01:10.98" />
                    <SPLIT distance="150" swimtime="00:01:48.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="443" swimtime="00:05:08.70" resultid="8265" heatid="10716" lane="0" entrytime="00:05:03.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                    <SPLIT distance="100" swimtime="00:01:11.76" />
                    <SPLIT distance="150" swimtime="00:01:50.36" />
                    <SPLIT distance="200" swimtime="00:02:30.03" />
                    <SPLIT distance="250" swimtime="00:03:10.22" />
                    <SPLIT distance="300" swimtime="00:03:50.82" />
                    <SPLIT distance="350" swimtime="00:04:30.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Magalhaes Dos Reis" birthdate="2010-05-05" gender="M" nation="BRA" license="356361" swrid="5600207" athleteid="8013" externalid="356361">
              <RESULTS>
                <RESULT eventid="1103" points="433" swimtime="00:00:29.43" resultid="8014" heatid="10506" lane="6" entrytime="00:00:30.22" entrycourse="LCM" />
                <RESULT eventid="1155" points="471" swimtime="00:00:59.62" resultid="8015" heatid="10549" lane="0" entrytime="00:00:59.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="457" swimtime="00:00:27.14" resultid="8016" heatid="10624" lane="4" entrytime="00:00:26.90" entrycourse="LCM" />
                <RESULT eventid="1219" points="362" swimtime="00:01:19.80" resultid="8017" heatid="10596" lane="8" entrytime="00:01:20.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="353" swimtime="00:02:41.20" resultid="8018" heatid="10650" lane="9" entrytime="00:02:36.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                    <SPLIT distance="100" swimtime="00:01:17.06" />
                    <SPLIT distance="150" swimtime="00:02:04.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="385" swimtime="00:02:20.14" resultid="8019" heatid="10662" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                    <SPLIT distance="100" swimtime="00:01:06.98" />
                    <SPLIT distance="150" swimtime="00:01:43.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Krupacz" birthdate="2008-04-18" gender="F" nation="BRA" license="329187" swrid="5634611" athleteid="7920" externalid="329187">
              <RESULTS>
                <RESULT eventid="1063" points="590" swimtime="00:02:26.77" resultid="7921" heatid="10473" lane="4" entrytime="00:02:26.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.87" />
                    <SPLIT distance="100" swimtime="00:01:10.42" />
                    <SPLIT distance="150" swimtime="00:01:48.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Albuquerque" birthdate="2012-08-17" gender="F" nation="BRA" license="369275" swrid="5602507" athleteid="8189" externalid="369275">
              <RESULTS>
                <RESULT eventid="1079" points="479" swimtime="00:02:55.70" resultid="8190" heatid="10485" lane="2" entrytime="00:02:58.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.09" />
                    <SPLIT distance="100" swimtime="00:01:24.10" />
                    <SPLIT distance="150" swimtime="00:02:10.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="340" swimtime="00:01:14.04" resultid="8191" heatid="10526" lane="2" entrytime="00:01:19.88" entrycourse="LCM" />
                <RESULT eventid="1227" points="367" swimtime="00:00:32.97" resultid="8192" heatid="10604" lane="2" entrytime="00:00:32.21" entrycourse="LCM" />
                <RESULT eventid="1211" points="522" swimtime="00:01:19.62" resultid="8193" heatid="10588" lane="4" entrytime="00:01:20.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="361" swimtime="00:02:57.09" resultid="8194" heatid="10641" lane="0" entrytime="00:03:02.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.80" />
                    <SPLIT distance="100" swimtime="00:01:31.00" />
                    <SPLIT distance="150" swimtime="00:02:16.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="264" swimtime="00:01:29.05" resultid="8195" heatid="10726" lane="4" entrytime="00:01:39.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Vieira Motta" birthdate="2009-09-19" gender="M" nation="BRA" license="339064" swrid="5600271" athleteid="7959" externalid="339064">
              <RESULTS>
                <RESULT eventid="1071" points="493" swimtime="00:02:21.58" resultid="7960" heatid="10480" lane="8" entrytime="00:02:19.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                    <SPLIT distance="100" swimtime="00:01:08.68" />
                    <SPLIT distance="150" swimtime="00:01:45.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="453" swimtime="00:01:00.41" resultid="7961" heatid="10548" lane="6" entrytime="00:01:00.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="486" swimtime="00:18:27.04" resultid="7962" heatid="10635" lane="1" entrytime="00:18:04.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                    <SPLIT distance="100" swimtime="00:01:07.24" />
                    <SPLIT distance="150" swimtime="00:01:43.13" />
                    <SPLIT distance="200" swimtime="00:02:19.27" />
                    <SPLIT distance="250" swimtime="00:02:55.75" />
                    <SPLIT distance="300" swimtime="00:03:32.36" />
                    <SPLIT distance="350" swimtime="00:04:08.78" />
                    <SPLIT distance="400" swimtime="00:04:45.82" />
                    <SPLIT distance="450" swimtime="00:05:22.66" />
                    <SPLIT distance="500" swimtime="00:05:59.85" />
                    <SPLIT distance="550" swimtime="00:06:36.93" />
                    <SPLIT distance="600" swimtime="00:07:14.57" />
                    <SPLIT distance="650" swimtime="00:07:52.15" />
                    <SPLIT distance="700" swimtime="00:08:29.51" />
                    <SPLIT distance="750" swimtime="00:09:06.92" />
                    <SPLIT distance="800" swimtime="00:09:44.48" />
                    <SPLIT distance="850" swimtime="00:10:21.45" />
                    <SPLIT distance="900" swimtime="00:10:59.17" />
                    <SPLIT distance="950" swimtime="00:11:36.72" />
                    <SPLIT distance="1000" swimtime="00:12:14.24" />
                    <SPLIT distance="1050" swimtime="00:12:51.49" />
                    <SPLIT distance="1100" swimtime="00:13:28.96" />
                    <SPLIT distance="1150" swimtime="00:14:05.93" />
                    <SPLIT distance="1200" swimtime="00:14:43.79" />
                    <SPLIT distance="1250" swimtime="00:15:21.19" />
                    <SPLIT distance="1300" swimtime="00:15:58.97" />
                    <SPLIT distance="1350" swimtime="00:16:36.06" />
                    <SPLIT distance="1400" swimtime="00:17:13.96" />
                    <SPLIT distance="1450" swimtime="00:17:50.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="478" swimtime="00:00:30.10" resultid="7963" heatid="10681" lane="2" />
                <RESULT eventid="1373" points="517" swimtime="00:01:04.29" resultid="7964" heatid="10742" lane="8" entrytime="00:01:03.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luisa" lastname="Della Villa Yang" birthdate="2012-10-08" gender="F" nation="BRA" license="369276" swrid="5588653" athleteid="8196" externalid="369276">
              <RESULTS>
                <RESULT eventid="1115" points="452" swimtime="00:19:58.68" resultid="8197" heatid="10511" lane="0" entrytime="00:20:11.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                    <SPLIT distance="100" swimtime="00:01:13.55" />
                    <SPLIT distance="150" swimtime="00:01:52.68" />
                    <SPLIT distance="200" swimtime="00:02:32.32" />
                    <SPLIT distance="250" swimtime="00:03:11.79" />
                    <SPLIT distance="300" swimtime="00:03:52.18" />
                    <SPLIT distance="350" swimtime="00:04:32.64" />
                    <SPLIT distance="400" swimtime="00:05:13.45" />
                    <SPLIT distance="450" swimtime="00:05:54.01" />
                    <SPLIT distance="500" swimtime="00:06:34.79" />
                    <SPLIT distance="550" swimtime="00:07:15.74" />
                    <SPLIT distance="600" swimtime="00:07:56.77" />
                    <SPLIT distance="650" swimtime="00:08:36.78" />
                    <SPLIT distance="700" swimtime="00:09:16.98" />
                    <SPLIT distance="750" swimtime="00:09:57.44" />
                    <SPLIT distance="800" swimtime="00:10:37.70" />
                    <SPLIT distance="850" swimtime="00:11:18.22" />
                    <SPLIT distance="900" swimtime="00:11:59.09" />
                    <SPLIT distance="950" swimtime="00:12:39.11" />
                    <SPLIT distance="1000" swimtime="00:13:19.33" />
                    <SPLIT distance="1050" swimtime="00:14:00.19" />
                    <SPLIT distance="1100" swimtime="00:14:40.33" />
                    <SPLIT distance="1150" swimtime="00:15:20.62" />
                    <SPLIT distance="1200" swimtime="00:16:01.15" />
                    <SPLIT distance="1250" swimtime="00:16:41.17" />
                    <SPLIT distance="1300" swimtime="00:17:21.47" />
                    <SPLIT distance="1350" swimtime="00:18:02.11" />
                    <SPLIT distance="1400" swimtime="00:18:41.82" />
                    <SPLIT distance="1450" swimtime="00:19:21.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="388" swimtime="00:06:02.31" resultid="8198" heatid="10519" lane="2" entrytime="00:06:11.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.13" />
                    <SPLIT distance="100" swimtime="00:01:29.67" />
                    <SPLIT distance="150" swimtime="00:02:16.90" />
                    <SPLIT distance="200" swimtime="00:03:02.89" />
                    <SPLIT distance="250" swimtime="00:03:55.17" />
                    <SPLIT distance="300" swimtime="00:04:47.03" />
                    <SPLIT distance="350" swimtime="00:05:25.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="482" swimtime="00:10:18.12" resultid="8199" heatid="10634" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="100" swimtime="00:01:12.59" />
                    <SPLIT distance="150" swimtime="00:01:51.41" />
                    <SPLIT distance="200" swimtime="00:02:29.80" />
                    <SPLIT distance="250" swimtime="00:03:08.55" />
                    <SPLIT distance="300" swimtime="00:03:47.29" />
                    <SPLIT distance="350" swimtime="00:04:26.61" />
                    <SPLIT distance="400" swimtime="00:05:06.49" />
                    <SPLIT distance="450" swimtime="00:05:46.11" />
                    <SPLIT distance="500" swimtime="00:06:25.66" />
                    <SPLIT distance="550" swimtime="00:07:05.06" />
                    <SPLIT distance="600" swimtime="00:07:44.23" />
                    <SPLIT distance="650" swimtime="00:08:23.28" />
                    <SPLIT distance="700" swimtime="00:09:02.28" />
                    <SPLIT distance="750" swimtime="00:09:40.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="404" swimtime="00:02:50.60" resultid="8200" heatid="10642" lane="9" entrytime="00:02:53.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                    <SPLIT distance="100" swimtime="00:01:21.31" />
                    <SPLIT distance="150" swimtime="00:02:13.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="479" swimtime="00:05:00.77" resultid="8201" heatid="10716" lane="1" entrytime="00:05:00.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                    <SPLIT distance="100" swimtime="00:01:09.40" />
                    <SPLIT distance="150" swimtime="00:01:47.16" />
                    <SPLIT distance="200" swimtime="00:02:25.77" />
                    <SPLIT distance="250" swimtime="00:03:04.77" />
                    <SPLIT distance="300" swimtime="00:03:43.85" />
                    <SPLIT distance="350" swimtime="00:04:22.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Leao" birthdate="2011-09-18" gender="M" nation="BRA" license="366880" swrid="5602553" athleteid="8034" externalid="366880">
              <RESULTS>
                <RESULT eventid="1123" points="430" swimtime="00:09:58.58" resultid="8035" heatid="10514" lane="8" entrytime="00:09:58.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                    <SPLIT distance="100" swimtime="00:01:10.57" />
                    <SPLIT distance="150" swimtime="00:01:48.10" />
                    <SPLIT distance="200" swimtime="00:02:25.45" />
                    <SPLIT distance="250" swimtime="00:03:03.58" />
                    <SPLIT distance="300" swimtime="00:03:41.28" />
                    <SPLIT distance="350" swimtime="00:04:19.71" />
                    <SPLIT distance="400" swimtime="00:04:57.60" />
                    <SPLIT distance="450" swimtime="00:05:36.01" />
                    <SPLIT distance="500" swimtime="00:06:14.11" />
                    <SPLIT distance="550" swimtime="00:06:52.59" />
                    <SPLIT distance="600" swimtime="00:07:30.94" />
                    <SPLIT distance="650" swimtime="00:08:08.83" />
                    <SPLIT distance="700" swimtime="00:08:46.30" />
                    <SPLIT distance="750" swimtime="00:09:23.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="431" swimtime="00:01:01.39" resultid="8036" heatid="10547" lane="8" entrytime="00:01:02.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="473" swimtime="00:18:36.86" resultid="8037" heatid="10636" lane="6" entrytime="00:19:05.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                    <SPLIT distance="100" swimtime="00:01:09.59" />
                    <SPLIT distance="150" swimtime="00:01:46.51" />
                    <SPLIT distance="200" swimtime="00:02:23.59" />
                    <SPLIT distance="250" swimtime="00:03:00.88" />
                    <SPLIT distance="300" swimtime="00:03:38.13" />
                    <SPLIT distance="350" swimtime="00:04:15.92" />
                    <SPLIT distance="400" swimtime="00:04:53.20" />
                    <SPLIT distance="450" swimtime="00:05:30.62" />
                    <SPLIT distance="500" swimtime="00:06:07.95" />
                    <SPLIT distance="550" swimtime="00:06:45.71" />
                    <SPLIT distance="600" swimtime="00:07:22.89" />
                    <SPLIT distance="650" swimtime="00:08:00.62" />
                    <SPLIT distance="700" swimtime="00:08:38.05" />
                    <SPLIT distance="750" swimtime="00:09:15.21" />
                    <SPLIT distance="800" swimtime="00:09:52.89" />
                    <SPLIT distance="850" swimtime="00:10:30.42" />
                    <SPLIT distance="900" swimtime="00:11:08.38" />
                    <SPLIT distance="950" swimtime="00:11:46.24" />
                    <SPLIT distance="1000" swimtime="00:12:24.06" />
                    <SPLIT distance="1050" swimtime="00:13:01.83" />
                    <SPLIT distance="1100" swimtime="00:13:39.42" />
                    <SPLIT distance="1150" swimtime="00:14:17.13" />
                    <SPLIT distance="1200" swimtime="00:14:55.01" />
                    <SPLIT distance="1250" swimtime="00:15:33.23" />
                    <SPLIT distance="1300" swimtime="00:16:11.04" />
                    <SPLIT distance="1350" swimtime="00:16:48.84" />
                    <SPLIT distance="1400" swimtime="00:17:26.38" />
                    <SPLIT distance="1450" swimtime="00:18:03.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="414" swimtime="00:00:28.05" resultid="8038" heatid="10619" lane="8" entrytime="00:00:29.95" entrycourse="LCM" />
                <RESULT eventid="1289" points="437" swimtime="00:02:14.38" resultid="8039" heatid="10670" lane="7" entrytime="00:02:16.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                    <SPLIT distance="100" swimtime="00:01:05.70" />
                    <SPLIT distance="150" swimtime="00:01:41.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="473" swimtime="00:04:42.36" resultid="8040" heatid="10722" lane="3" entrytime="00:04:43.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.34" />
                    <SPLIT distance="100" swimtime="00:01:06.65" />
                    <SPLIT distance="150" swimtime="00:01:42.80" />
                    <SPLIT distance="200" swimtime="00:02:19.38" />
                    <SPLIT distance="250" swimtime="00:02:56.04" />
                    <SPLIT distance="300" swimtime="00:03:33.22" />
                    <SPLIT distance="350" swimtime="00:04:09.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Spadari Soso" birthdate="2012-12-28" gender="F" nation="BRA" license="377313" swrid="5588921" athleteid="8353" externalid="377313">
              <RESULTS>
                <RESULT eventid="1079" points="394" swimtime="00:03:07.62" resultid="8354" heatid="10483" lane="4" entrytime="00:03:08.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.23" />
                    <SPLIT distance="100" swimtime="00:01:29.68" />
                    <SPLIT distance="150" swimtime="00:02:18.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="486" swimtime="00:01:05.77" resultid="8355" heatid="10532" lane="7" entrytime="00:01:05.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="442" swimtime="00:00:30.98" resultid="8356" heatid="10606" lane="2" entrytime="00:00:30.96" entrycourse="LCM" />
                <RESULT eventid="1211" points="365" swimtime="00:01:29.72" resultid="8357" heatid="10586" lane="4" entrytime="00:01:27.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="498" swimtime="00:02:21.58" resultid="8358" heatid="10657" lane="4" entrytime="00:02:28.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.84" />
                    <SPLIT distance="100" swimtime="00:01:09.68" />
                    <SPLIT distance="150" swimtime="00:01:46.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="440" swimtime="00:05:09.44" resultid="8359" heatid="10714" lane="3" entrytime="00:05:16.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.12" />
                    <SPLIT distance="100" swimtime="00:01:14.69" />
                    <SPLIT distance="150" swimtime="00:01:54.98" />
                    <SPLIT distance="200" swimtime="00:02:35.86" />
                    <SPLIT distance="250" swimtime="00:03:15.52" />
                    <SPLIT distance="300" swimtime="00:03:54.91" />
                    <SPLIT distance="350" swimtime="00:04:32.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Carneiro Silva" birthdate="2011-02-21" gender="F" nation="BRA" license="390924" swrid="5602522" athleteid="8323" externalid="390924">
              <RESULTS>
                <RESULT eventid="1063" points="420" swimtime="00:02:44.35" resultid="8324" heatid="10472" lane="4" entrytime="00:02:44.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                    <SPLIT distance="100" swimtime="00:01:16.68" />
                    <SPLIT distance="150" swimtime="00:02:00.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="434" swimtime="00:01:08.28" resultid="8325" heatid="10530" lane="4" entrytime="00:01:08.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="449" swimtime="00:00:30.83" resultid="8326" heatid="10606" lane="8" entrytime="00:00:31.15" entrycourse="LCM" />
                <RESULT eventid="1265" points="385" swimtime="00:02:53.32" resultid="8327" heatid="10641" lane="1" entrytime="00:03:01.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.32" />
                    <SPLIT distance="100" swimtime="00:01:21.63" />
                    <SPLIT distance="150" swimtime="00:02:15.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="362" swimtime="00:02:37.42" resultid="8328" heatid="10657" lane="0" entrytime="00:02:30.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                    <SPLIT distance="100" swimtime="00:01:15.23" />
                    <SPLIT distance="150" swimtime="00:01:56.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="422" swimtime="00:01:16.16" resultid="8329" heatid="10731" lane="3" entrytime="00:01:16.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maryna" lastname="Monegat Fachin" birthdate="2008-01-02" gender="F" nation="BRA" license="341528" swrid="5634727" athleteid="8399" externalid="341528">
              <RESULTS>
                <RESULT eventid="1115" points="635" swimtime="00:17:50.82" resultid="8400" heatid="10511" lane="3" entrytime="00:18:17.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                    <SPLIT distance="100" swimtime="00:01:08.32" />
                    <SPLIT distance="150" swimtime="00:01:43.67" />
                    <SPLIT distance="200" swimtime="00:02:19.05" />
                    <SPLIT distance="250" swimtime="00:02:54.84" />
                    <SPLIT distance="300" swimtime="00:03:30.63" />
                    <SPLIT distance="350" swimtime="00:04:06.46" />
                    <SPLIT distance="400" swimtime="00:04:41.62" />
                    <SPLIT distance="450" swimtime="00:05:17.11" />
                    <SPLIT distance="500" swimtime="00:05:52.42" />
                    <SPLIT distance="550" swimtime="00:06:27.95" />
                    <SPLIT distance="600" swimtime="00:07:03.14" />
                    <SPLIT distance="650" swimtime="00:07:39.10" />
                    <SPLIT distance="700" swimtime="00:08:14.79" />
                    <SPLIT distance="750" swimtime="00:08:50.63" />
                    <SPLIT distance="800" swimtime="00:09:26.31" />
                    <SPLIT distance="850" swimtime="00:10:02.66" />
                    <SPLIT distance="900" swimtime="00:10:38.75" />
                    <SPLIT distance="950" swimtime="00:11:14.85" />
                    <SPLIT distance="1000" swimtime="00:11:50.57" />
                    <SPLIT distance="1050" swimtime="00:12:26.68" />
                    <SPLIT distance="1100" swimtime="00:13:02.71" />
                    <SPLIT distance="1150" swimtime="00:13:38.67" />
                    <SPLIT distance="1200" swimtime="00:14:14.67" />
                    <SPLIT distance="1250" swimtime="00:14:51.01" />
                    <SPLIT distance="1300" swimtime="00:15:27.08" />
                    <SPLIT distance="1350" swimtime="00:16:03.38" />
                    <SPLIT distance="1400" swimtime="00:16:39.96" />
                    <SPLIT distance="1450" swimtime="00:17:16.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Vitoria Kuzmann Cercal" birthdate="2009-04-10" gender="F" nation="BRA" license="339082" swrid="5600274" athleteid="7949" externalid="339082">
              <RESULTS>
                <RESULT eventid="1095" points="431" swimtime="00:00:32.32" resultid="7950" heatid="10494" lane="1" />
                <RESULT eventid="1147" points="545" swimtime="00:01:03.27" resultid="7951" heatid="10534" lane="0" entrytime="00:01:03.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="510" swimtime="00:00:29.54" resultid="7952" heatid="10608" lane="4" entrytime="00:00:29.27" entrycourse="LCM" />
                <RESULT eventid="1281" points="455" swimtime="00:02:25.88" resultid="7953" heatid="10657" lane="3" entrytime="00:02:28.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                    <SPLIT distance="100" swimtime="00:01:09.64" />
                    <SPLIT distance="150" swimtime="00:01:47.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Fernandes  Dos Reis" birthdate="2012-09-18" gender="M" nation="BRA" license="369279" swrid="5588696" athleteid="8215" externalid="369279">
              <RESULTS>
                <RESULT eventid="1103" points="289" swimtime="00:00:33.68" resultid="8216" heatid="10504" lane="7" entrytime="00:00:33.97" entrycourse="LCM" />
                <RESULT eventid="1171" points="245" swimtime="00:02:56.26" resultid="8217" heatid="10556" lane="1" entrytime="00:02:55.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                    <SPLIT distance="100" swimtime="00:01:21.40" />
                    <SPLIT distance="150" swimtime="00:02:09.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" status="DNS" swimtime="00:00:00.00" resultid="8218" heatid="10616" lane="5" entrytime="00:00:31.73" entrycourse="LCM" />
                <RESULT eventid="1273" points="293" swimtime="00:02:51.45" resultid="8219" heatid="10647" lane="3" entrytime="00:02:55.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.49" />
                    <SPLIT distance="100" swimtime="00:01:23.15" />
                    <SPLIT distance="150" swimtime="00:02:16.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="279" swimtime="00:01:15.61" resultid="8220" heatid="10706" lane="4" entrytime="00:01:16.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Trevisan" birthdate="2000-11-28" gender="M" nation="BRA" license="346847" swrid="5600266" athleteid="8305" externalid="346847">
              <RESULTS>
                <RESULT eventid="1235" points="607" swimtime="00:00:24.69" resultid="8306" heatid="10628" lane="2" entrytime="00:00:24.39" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Pedro Pasqual" birthdate="2009-06-17" gender="M" nation="BRA" license="386136" swrid="5600232" athleteid="7908" externalid="386136">
              <RESULTS>
                <RESULT eventid="1071" status="DNS" swimtime="00:00:00.00" resultid="7909" heatid="10480" lane="6" entrytime="00:02:14.97" entrycourse="LCM" />
                <RESULT eventid="1155" points="599" swimtime="00:00:55.02" resultid="7910" heatid="10551" lane="6" entrytime="00:00:55.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="547" swimtime="00:02:04.65" resultid="7911" heatid="10672" lane="0" entrytime="00:02:09.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.78" />
                    <SPLIT distance="100" swimtime="00:01:00.17" />
                    <SPLIT distance="150" swimtime="00:01:34.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="630" swimtime="00:01:00.19" resultid="7912" heatid="10742" lane="5" entrytime="00:01:00.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Muxfeldt" birthdate="2011-05-13" gender="F" nation="BRA" license="366903" swrid="5602563" athleteid="8076" externalid="366903">
              <RESULTS>
                <RESULT eventid="1115" points="438" swimtime="00:20:11.67" resultid="8077" heatid="10512" lane="4" entrytime="00:20:22.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                    <SPLIT distance="100" swimtime="00:01:15.96" />
                    <SPLIT distance="150" swimtime="00:01:55.41" />
                    <SPLIT distance="200" swimtime="00:02:35.86" />
                    <SPLIT distance="250" swimtime="00:03:17.43" />
                    <SPLIT distance="300" swimtime="00:03:58.59" />
                    <SPLIT distance="350" swimtime="00:04:38.69" />
                    <SPLIT distance="400" swimtime="00:05:19.36" />
                    <SPLIT distance="450" swimtime="00:06:00.65" />
                    <SPLIT distance="500" swimtime="00:06:41.71" />
                    <SPLIT distance="550" swimtime="00:07:22.21" />
                    <SPLIT distance="600" swimtime="00:08:02.94" />
                    <SPLIT distance="650" swimtime="00:08:43.27" />
                    <SPLIT distance="700" swimtime="00:09:24.41" />
                    <SPLIT distance="750" swimtime="00:10:05.27" />
                    <SPLIT distance="800" swimtime="00:10:45.59" />
                    <SPLIT distance="850" swimtime="00:11:25.26" />
                    <SPLIT distance="900" swimtime="00:12:06.37" />
                    <SPLIT distance="950" swimtime="00:12:47.61" />
                    <SPLIT distance="1000" swimtime="00:13:28.34" />
                    <SPLIT distance="1050" swimtime="00:14:08.96" />
                    <SPLIT distance="1100" swimtime="00:14:49.63" />
                    <SPLIT distance="1150" swimtime="00:15:30.84" />
                    <SPLIT distance="1200" swimtime="00:16:11.42" />
                    <SPLIT distance="1250" swimtime="00:16:52.04" />
                    <SPLIT distance="1300" swimtime="00:17:32.91" />
                    <SPLIT distance="1350" swimtime="00:18:13.50" />
                    <SPLIT distance="1400" swimtime="00:18:54.76" />
                    <SPLIT distance="1450" swimtime="00:19:34.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="347" swimtime="00:03:15.69" resultid="8078" heatid="10484" lane="3" entrytime="00:03:04.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.41" />
                    <SPLIT distance="100" swimtime="00:01:33.92" />
                    <SPLIT distance="150" swimtime="00:02:26.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="483" swimtime="00:01:05.87" resultid="8079" heatid="10531" lane="0" entrytime="00:01:07.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="444" swimtime="00:00:30.93" resultid="8080" heatid="10606" lane="6" entrytime="00:00:30.86" entrycourse="LCM" />
                <RESULT eventid="1211" points="345" swimtime="00:01:31.35" resultid="8081" heatid="10587" lane="6" entrytime="00:01:25.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="509" swimtime="00:02:20.48" resultid="8082" heatid="10658" lane="6" entrytime="00:02:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.88" />
                    <SPLIT distance="100" swimtime="00:01:09.33" />
                    <SPLIT distance="150" swimtime="00:01:45.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Clara Fernandes Pereira" birthdate="2009-11-19" gender="F" nation="BRA" license="344340" swrid="5600137" athleteid="7821" externalid="344340">
              <RESULTS>
                <RESULT eventid="1079" points="445" swimtime="00:03:00.09" resultid="7822" heatid="10485" lane="9" entrytime="00:03:02.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.16" />
                    <SPLIT distance="100" swimtime="00:01:26.81" />
                    <SPLIT distance="150" swimtime="00:02:14.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="437" swimtime="00:01:24.50" resultid="7823" heatid="10583" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="540" swimtime="00:02:17.74" resultid="7824" heatid="10660" lane="6" entrytime="00:02:17.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                    <SPLIT distance="100" swimtime="00:01:06.38" />
                    <SPLIT distance="150" swimtime="00:01:41.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="517" swimtime="00:04:53.26" resultid="7825" heatid="10716" lane="5" entrytime="00:04:47.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.26" />
                    <SPLIT distance="100" swimtime="00:01:09.33" />
                    <SPLIT distance="150" swimtime="00:01:46.04" />
                    <SPLIT distance="200" swimtime="00:02:23.37" />
                    <SPLIT distance="250" swimtime="00:03:00.70" />
                    <SPLIT distance="300" swimtime="00:03:38.24" />
                    <SPLIT distance="350" swimtime="00:04:15.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tiago" lastname="Lacerda" birthdate="2011-05-09" gender="M" nation="BRA" license="366909" swrid="5602550" athleteid="8111" externalid="366909">
              <RESULTS>
                <RESULT eventid="1071" points="370" swimtime="00:02:35.82" resultid="8112" heatid="10475" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                    <SPLIT distance="100" swimtime="00:01:15.61" />
                    <SPLIT distance="150" swimtime="00:01:56.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="398" swimtime="00:05:29.58" resultid="8113" heatid="10522" lane="8" entrytime="00:05:35.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                    <SPLIT distance="100" swimtime="00:01:16.97" />
                    <SPLIT distance="150" swimtime="00:01:59.54" />
                    <SPLIT distance="200" swimtime="00:02:40.04" />
                    <SPLIT distance="250" swimtime="00:03:28.16" />
                    <SPLIT distance="300" swimtime="00:04:14.93" />
                    <SPLIT distance="350" swimtime="00:04:53.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="305" swimtime="00:01:24.50" resultid="8114" heatid="10594" lane="1" entrytime="00:01:27.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="417" swimtime="00:02:32.50" resultid="8115" heatid="10650" lane="6" entrytime="00:02:31.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                    <SPLIT distance="100" swimtime="00:01:13.56" />
                    <SPLIT distance="150" swimtime="00:01:58.77" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 9:12)" eventid="1341" status="DSQ" swimtime="00:01:11.17" resultid="8116" heatid="10704" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="380" swimtime="00:01:11.20" resultid="8117" heatid="10739" lane="8" entrytime="00:01:11.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rene" lastname="Osternack Erbe" birthdate="2011-04-03" gender="M" nation="BRA" license="366907" swrid="5588842" athleteid="8097" externalid="366907">
              <RESULTS>
                <RESULT eventid="1103" points="276" swimtime="00:00:34.17" resultid="8098" heatid="10500" lane="3" />
                <RESULT eventid="1071" points="346" swimtime="00:02:39.35" resultid="8099" heatid="10477" lane="1" entrytime="00:02:42.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                    <SPLIT distance="100" swimtime="00:01:17.89" />
                    <SPLIT distance="150" swimtime="00:01:59.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="328" swimtime="00:01:07.25" resultid="8100" heatid="10542" lane="6" entrytime="00:01:09.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="317" swimtime="00:00:30.66" resultid="8101" heatid="10618" lane="0" entrytime="00:00:30.89" entrycourse="LCM" />
                <RESULT eventid="1305" points="319" swimtime="00:00:34.45" resultid="8102" heatid="10684" lane="4" entrytime="00:00:36.68" entrycourse="LCM" />
                <RESULT eventid="1373" points="346" swimtime="00:01:13.45" resultid="8103" heatid="10738" lane="3" entrytime="00:01:14.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Giuseppe Bulla Lanaro" birthdate="2007-05-22" gender="M" nation="BRA" license="331630" swrid="5600174" athleteid="7892" externalid="331630">
              <RESULTS>
                <RESULT eventid="1123" points="558" swimtime="00:09:09.05" resultid="7893" heatid="10513" lane="4" entrytime="00:08:51.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                    <SPLIT distance="100" swimtime="00:01:02.47" />
                    <SPLIT distance="150" swimtime="00:01:36.14" />
                    <SPLIT distance="200" swimtime="00:02:10.26" />
                    <SPLIT distance="250" swimtime="00:02:43.95" />
                    <SPLIT distance="300" swimtime="00:03:17.86" />
                    <SPLIT distance="350" swimtime="00:03:52.02" />
                    <SPLIT distance="400" swimtime="00:04:26.37" />
                    <SPLIT distance="450" swimtime="00:05:00.68" />
                    <SPLIT distance="500" swimtime="00:05:35.28" />
                    <SPLIT distance="550" swimtime="00:06:10.37" />
                    <SPLIT distance="600" swimtime="00:06:46.44" />
                    <SPLIT distance="650" swimtime="00:07:22.83" />
                    <SPLIT distance="700" swimtime="00:07:59.53" />
                    <SPLIT distance="750" swimtime="00:08:35.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="628" swimtime="00:00:54.17" resultid="7894" heatid="10552" lane="1" entrytime="00:00:53.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="549" swimtime="00:00:25.53" resultid="7895" heatid="10627" lane="2" entrytime="00:00:25.22" entrycourse="LCM" />
                <RESULT eventid="1289" points="651" swimtime="00:01:57.65" resultid="7896" heatid="10674" lane="2" entrytime="00:01:57.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.83" />
                    <SPLIT distance="100" swimtime="00:00:57.66" />
                    <SPLIT distance="150" swimtime="00:01:27.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="651" swimtime="00:04:13.88" resultid="7897" heatid="10724" lane="5" entrytime="00:04:12.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.69" />
                    <SPLIT distance="100" swimtime="00:01:00.09" />
                    <SPLIT distance="150" swimtime="00:01:31.99" />
                    <SPLIT distance="200" swimtime="00:02:04.25" />
                    <SPLIT distance="250" swimtime="00:02:36.36" />
                    <SPLIT distance="300" swimtime="00:03:08.76" />
                    <SPLIT distance="350" swimtime="00:03:41.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martina" lastname="Mayer Paludetto" birthdate="2012-10-30" gender="F" nation="BRA" license="369264" swrid="5588811" athleteid="8149" externalid="369264">
              <RESULTS>
                <RESULT eventid="1063" points="409" swimtime="00:02:45.80" resultid="8150" heatid="10472" lane="8" entrytime="00:02:48.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                    <SPLIT distance="100" swimtime="00:01:18.79" />
                    <SPLIT distance="150" swimtime="00:02:03.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="572" swimtime="00:01:02.26" resultid="8151" heatid="10531" lane="3" entrytime="00:01:06.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="508" swimtime="00:10:07.18" resultid="8152" heatid="10634" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                    <SPLIT distance="100" swimtime="00:01:07.51" />
                    <SPLIT distance="150" swimtime="00:01:45.24" />
                    <SPLIT distance="200" swimtime="00:02:24.11" />
                    <SPLIT distance="250" swimtime="00:03:03.03" />
                    <SPLIT distance="300" swimtime="00:03:42.11" />
                    <SPLIT distance="350" swimtime="00:04:20.99" />
                    <SPLIT distance="400" swimtime="00:04:59.98" />
                    <SPLIT distance="450" swimtime="00:05:38.99" />
                    <SPLIT distance="500" swimtime="00:06:18.32" />
                    <SPLIT distance="550" swimtime="00:06:57.72" />
                    <SPLIT distance="600" swimtime="00:07:37.09" />
                    <SPLIT distance="650" swimtime="00:08:16.05" />
                    <SPLIT distance="700" swimtime="00:08:54.00" />
                    <SPLIT distance="750" swimtime="00:09:30.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="532" swimtime="00:02:18.46" resultid="8153" heatid="10660" lane="1" entrytime="00:02:18.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.20" />
                    <SPLIT distance="100" swimtime="00:01:05.76" />
                    <SPLIT distance="150" swimtime="00:01:42.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="546" swimtime="00:04:47.92" resultid="8154" heatid="10716" lane="3" entrytime="00:04:53.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                    <SPLIT distance="100" swimtime="00:01:08.11" />
                    <SPLIT distance="150" swimtime="00:01:43.82" />
                    <SPLIT distance="200" swimtime="00:02:21.50" />
                    <SPLIT distance="250" swimtime="00:02:58.29" />
                    <SPLIT distance="300" swimtime="00:03:35.68" />
                    <SPLIT distance="350" swimtime="00:04:12.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="398" swimtime="00:01:17.61" resultid="8155" heatid="10730" lane="8" entrytime="00:01:19.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Szpak De Vasconcelos" birthdate="2012-06-29" gender="M" nation="BRA" license="369271" swrid="5588928" athleteid="8176" externalid="369271">
              <RESULTS>
                <RESULT eventid="1087" points="338" swimtime="00:02:59.98" resultid="8177" heatid="10489" lane="4" entrytime="00:03:01.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.90" />
                    <SPLIT distance="100" swimtime="00:01:27.36" />
                    <SPLIT distance="150" swimtime="00:02:14.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="357" swimtime="00:01:05.36" resultid="8178" heatid="10544" lane="9" entrytime="00:01:06.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="331" swimtime="00:01:22.22" resultid="8179" heatid="10595" lane="2" entrytime="00:01:22.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="323" swimtime="00:02:28.52" resultid="8180" heatid="10667" lane="1" entrytime="00:02:30.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                    <SPLIT distance="100" swimtime="00:01:10.72" />
                    <SPLIT distance="150" swimtime="00:01:49.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="282" swimtime="00:01:18.65" resultid="8181" heatid="10736" lane="5" entrytime="00:01:20.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietra" lastname="Ruschel Carvalho" birthdate="2009-03-21" gender="F" nation="BRA" license="324999" swrid="5600250" athleteid="7826" externalid="324999">
              <RESULTS>
                <RESULT eventid="1095" points="508" swimtime="00:00:30.60" resultid="7827" heatid="10498" lane="7" entrytime="00:00:31.57" entrycourse="LCM" />
                <RESULT eventid="1147" points="647" swimtime="00:00:59.78" resultid="7828" heatid="10534" lane="4" entrytime="00:00:59.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="648" swimtime="00:00:27.28" resultid="7829" heatid="10609" lane="4" entrytime="00:00:26.92" entrycourse="LCM" />
                <RESULT eventid="1281" points="560" swimtime="00:02:16.14" resultid="7830" heatid="10660" lane="3" entrytime="00:02:11.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                    <SPLIT distance="100" swimtime="00:01:03.34" />
                    <SPLIT distance="150" swimtime="00:01:39.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="438" swimtime="00:01:12.61" resultid="7831" heatid="10699" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Prosdocimo" birthdate="2010-11-23" gender="F" nation="BRA" license="356251" swrid="5600238" athleteid="7985" externalid="356251">
              <RESULTS>
                <RESULT eventid="1115" points="396" swimtime="00:20:52.84" resultid="7986" heatid="10511" lane="9" entrytime="00:20:18.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                    <SPLIT distance="100" swimtime="00:01:18.23" />
                    <SPLIT distance="150" swimtime="00:01:59.35" />
                    <SPLIT distance="200" swimtime="00:02:41.36" />
                    <SPLIT distance="250" swimtime="00:03:23.02" />
                    <SPLIT distance="300" swimtime="00:04:05.26" />
                    <SPLIT distance="350" swimtime="00:04:47.51" />
                    <SPLIT distance="400" swimtime="00:05:30.27" />
                    <SPLIT distance="450" swimtime="00:06:12.62" />
                    <SPLIT distance="500" swimtime="00:06:55.26" />
                    <SPLIT distance="550" swimtime="00:07:37.97" />
                    <SPLIT distance="600" swimtime="00:08:21.18" />
                    <SPLIT distance="650" swimtime="00:09:03.85" />
                    <SPLIT distance="700" swimtime="00:09:46.67" />
                    <SPLIT distance="750" swimtime="00:10:29.03" />
                    <SPLIT distance="800" swimtime="00:11:11.52" />
                    <SPLIT distance="850" swimtime="00:11:53.03" />
                    <SPLIT distance="900" swimtime="00:12:34.50" />
                    <SPLIT distance="950" swimtime="00:13:16.50" />
                    <SPLIT distance="1000" swimtime="00:13:58.22" />
                    <SPLIT distance="1050" swimtime="00:14:40.40" />
                    <SPLIT distance="1100" swimtime="00:15:22.63" />
                    <SPLIT distance="1150" swimtime="00:16:04.53" />
                    <SPLIT distance="1200" swimtime="00:16:46.72" />
                    <SPLIT distance="1250" swimtime="00:17:28.44" />
                    <SPLIT distance="1300" swimtime="00:18:09.37" />
                    <SPLIT distance="1350" swimtime="00:18:51.05" />
                    <SPLIT distance="1400" swimtime="00:19:32.74" />
                    <SPLIT distance="1450" swimtime="00:20:13.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="381" swimtime="00:02:49.82" resultid="7987" heatid="10472" lane="2" entrytime="00:02:46.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                    <SPLIT distance="100" swimtime="00:01:23.46" />
                    <SPLIT distance="150" swimtime="00:02:06.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="478" swimtime="00:01:06.10" resultid="7988" heatid="10533" lane="9" entrytime="00:01:05.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="469" swimtime="00:00:30.38" resultid="7989" heatid="10607" lane="1" entrytime="00:00:30.46" entrycourse="LCM" />
                <RESULT eventid="1265" points="362" swimtime="00:02:56.92" resultid="7990" heatid="10639" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                    <SPLIT distance="100" swimtime="00:01:22.94" />
                    <SPLIT distance="150" swimtime="00:02:21.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="389" swimtime="00:01:18.25" resultid="7991" heatid="10731" lane="5" entrytime="00:01:15.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olivia" lastname="Jeger" birthdate="2004-12-19" gender="F" nation="BRA" license="325493" swrid="5600193" athleteid="8321" externalid="325493" level="UNIDOMBOSC">
              <RESULTS>
                <RESULT eventid="1115" points="642" swimtime="00:17:46.56" resultid="8322" heatid="10511" lane="5" entrytime="00:17:57.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.42" />
                    <SPLIT distance="100" swimtime="00:01:07.35" />
                    <SPLIT distance="150" swimtime="00:01:42.59" />
                    <SPLIT distance="200" swimtime="00:02:18.22" />
                    <SPLIT distance="250" swimtime="00:02:53.63" />
                    <SPLIT distance="300" swimtime="00:03:29.62" />
                    <SPLIT distance="350" swimtime="00:04:05.11" />
                    <SPLIT distance="400" swimtime="00:04:41.10" />
                    <SPLIT distance="450" swimtime="00:05:16.58" />
                    <SPLIT distance="500" swimtime="00:05:52.55" />
                    <SPLIT distance="550" swimtime="00:06:28.14" />
                    <SPLIT distance="600" swimtime="00:07:04.15" />
                    <SPLIT distance="650" swimtime="00:07:39.69" />
                    <SPLIT distance="700" swimtime="00:08:15.76" />
                    <SPLIT distance="750" swimtime="00:08:51.39" />
                    <SPLIT distance="800" swimtime="00:09:27.69" />
                    <SPLIT distance="850" swimtime="00:10:03.37" />
                    <SPLIT distance="900" swimtime="00:10:39.53" />
                    <SPLIT distance="950" swimtime="00:11:15.06" />
                    <SPLIT distance="1000" swimtime="00:11:51.06" />
                    <SPLIT distance="1050" swimtime="00:12:26.70" />
                    <SPLIT distance="1100" swimtime="00:13:02.80" />
                    <SPLIT distance="1150" swimtime="00:13:38.40" />
                    <SPLIT distance="1200" swimtime="00:14:14.78" />
                    <SPLIT distance="1250" swimtime="00:14:49.91" />
                    <SPLIT distance="1300" swimtime="00:15:25.94" />
                    <SPLIT distance="1350" swimtime="00:16:01.17" />
                    <SPLIT distance="1400" swimtime="00:16:37.02" />
                    <SPLIT distance="1450" swimtime="00:17:12.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Vanzo Assumpcao" birthdate="2012-05-15" gender="M" nation="BRA" license="369258" swrid="5588942" athleteid="8122" externalid="369258">
              <RESULTS>
                <RESULT eventid="1071" status="DNS" swimtime="00:00:00.00" resultid="8123" heatid="10475" lane="9" />
                <RESULT eventid="1171" status="DNS" swimtime="00:00:00.00" resultid="8124" heatid="10556" lane="4" entrytime="00:02:40.71" entrycourse="LCM" />
                <RESULT eventid="1235" status="DNS" swimtime="00:00:00.00" resultid="8125" heatid="10611" lane="3" />
                <RESULT eventid="1289" points="429" swimtime="00:02:15.14" resultid="8126" heatid="10670" lane="0" entrytime="00:02:18.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.81" />
                    <SPLIT distance="100" swimtime="00:01:06.83" />
                    <SPLIT distance="150" swimtime="00:01:41.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="404" swimtime="00:01:06.87" resultid="8127" heatid="10709" lane="9" entrytime="00:01:07.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="376" swimtime="00:01:11.49" resultid="8128" heatid="10738" lane="2" entrytime="00:01:14.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Novak Bredt" birthdate="2009-09-08" gender="F" nation="BRA" license="338909" swrid="5622297" athleteid="7878" externalid="338909">
              <RESULTS>
                <RESULT eventid="1079" points="475" swimtime="00:02:56.24" resultid="7879" heatid="10485" lane="4" entrytime="00:02:56.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.97" />
                    <SPLIT distance="100" swimtime="00:01:23.47" />
                    <SPLIT distance="150" swimtime="00:02:10.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="489" swimtime="00:00:37.01" resultid="7880" heatid="10564" lane="2" entrytime="00:00:38.16" entrycourse="LCM" />
                <RESULT eventid="1211" points="497" swimtime="00:01:20.96" resultid="7881" heatid="10588" lane="6" entrytime="00:01:21.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="463" swimtime="00:02:42.92" resultid="7882" heatid="10644" lane="9" entrytime="00:02:42.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.73" />
                    <SPLIT distance="100" swimtime="00:01:16.40" />
                    <SPLIT distance="150" swimtime="00:02:03.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="400" swimtime="00:01:14.83" resultid="7883" heatid="10701" lane="5" entrytime="00:01:16.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Brandt De Macedo" birthdate="2006-04-22" gender="M" nation="BRA" license="296648" swrid="5622265" athleteid="7857" externalid="296648">
              <RESULTS>
                <RESULT eventid="1357" points="759" swimtime="00:04:01.19" resultid="7858" heatid="10724" lane="4" entrytime="00:04:04.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.14" />
                    <SPLIT distance="100" swimtime="00:00:58.27" />
                    <SPLIT distance="150" swimtime="00:01:28.57" />
                    <SPLIT distance="200" swimtime="00:01:59.29" />
                    <SPLIT distance="250" swimtime="00:02:29.96" />
                    <SPLIT distance="300" swimtime="00:03:01.04" />
                    <SPLIT distance="350" swimtime="00:03:31.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio" lastname="Sabedotti" birthdate="2002-07-07" gender="M" nation="BRA" license="134704" swrid="5600252" athleteid="7969" externalid="134704" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1219" points="661" swimtime="00:01:05.27" resultid="7970" heatid="10599" lane="2" entrytime="00:01:04.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Moreira Segadaes" birthdate="2008-05-15" gender="M" nation="BRA" license="331574" swrid="5600220" athleteid="7851" externalid="331574">
              <RESULTS>
                <RESULT eventid="1187" points="586" swimtime="00:00:31.00" resultid="7852" heatid="10575" lane="1" entrytime="00:00:30.89" entrycourse="LCM" />
                <RESULT eventid="1235" points="498" swimtime="00:00:26.37" resultid="7853" heatid="10611" lane="7" />
                <RESULT eventid="1219" points="576" swimtime="00:01:08.33" resultid="7854" heatid="10599" lane="8" entrytime="00:01:07.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruna" lastname="Bussmann" birthdate="2007-01-16" gender="F" nation="BRA" license="313781" swrid="5579983" athleteid="7855" externalid="313781">
              <RESULTS>
                <RESULT eventid="1211" points="598" swimtime="00:01:16.11" resultid="7856" heatid="10589" lane="4" entrytime="00:01:14.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gael" lastname="Gluck" birthdate="2011-01-28" gender="M" nation="BRA" license="366891" swrid="5588726" athleteid="8048" externalid="366891">
              <RESULTS>
                <RESULT eventid="1087" points="411" swimtime="00:02:48.64" resultid="8049" heatid="10491" lane="8" entrytime="00:02:48.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.42" />
                    <SPLIT distance="100" swimtime="00:01:19.54" />
                    <SPLIT distance="150" swimtime="00:02:03.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="465" swimtime="00:00:59.86" resultid="8050" heatid="10546" lane="2" entrytime="00:01:02.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="402" swimtime="00:00:28.33" resultid="8051" heatid="10621" lane="4" entrytime="00:00:28.33" entrycourse="LCM" />
                <RESULT eventid="1219" points="369" swimtime="00:01:19.27" resultid="8052" heatid="10597" lane="0" entrytime="00:01:18.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="506" swimtime="00:02:07.96" resultid="8053" heatid="10671" lane="5" entrytime="00:02:11.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.20" />
                    <SPLIT distance="100" swimtime="00:01:02.26" />
                    <SPLIT distance="150" swimtime="00:01:34.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="510" swimtime="00:04:35.35" resultid="8054" heatid="10723" lane="9" entrytime="00:04:39.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                    <SPLIT distance="100" swimtime="00:01:05.92" />
                    <SPLIT distance="150" swimtime="00:01:40.73" />
                    <SPLIT distance="200" swimtime="00:02:15.97" />
                    <SPLIT distance="250" swimtime="00:02:51.01" />
                    <SPLIT distance="300" swimtime="00:03:26.06" />
                    <SPLIT distance="350" swimtime="00:04:01.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="LIV" lastname="Carvalho" birthdate="2011-09-13" gender="F" nation="BRA" license="366899" swrid="5602524" athleteid="8069" externalid="366899">
              <RESULTS>
                <RESULT eventid="1079" points="397" swimtime="00:03:07.02" resultid="8070" heatid="10484" lane="7" entrytime="00:03:06.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.77" />
                    <SPLIT distance="100" swimtime="00:01:30.28" />
                    <SPLIT distance="150" swimtime="00:02:19.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="333" swimtime="00:00:42.07" resultid="8071" heatid="10563" lane="6" entrytime="00:00:40.85" entrycourse="LCM" />
                <RESULT eventid="1147" points="358" swimtime="00:01:12.77" resultid="8072" heatid="10527" lane="3" entrytime="00:01:15.19" entrycourse="LCM" />
                <RESULT eventid="1249" points="355" swimtime="00:11:24.50" resultid="8073" heatid="10633" lane="2" entrytime="00:11:35.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                    <SPLIT distance="100" swimtime="00:01:18.75" />
                    <SPLIT distance="150" swimtime="00:01:59.76" />
                    <SPLIT distance="200" swimtime="00:02:42.33" />
                    <SPLIT distance="250" swimtime="00:03:25.34" />
                    <SPLIT distance="300" swimtime="00:04:09.68" />
                    <SPLIT distance="350" swimtime="00:04:53.24" />
                    <SPLIT distance="400" swimtime="00:05:37.77" />
                    <SPLIT distance="450" swimtime="00:06:20.48" />
                    <SPLIT distance="500" swimtime="00:07:04.56" />
                    <SPLIT distance="550" swimtime="00:07:48.31" />
                    <SPLIT distance="600" swimtime="00:08:32.69" />
                    <SPLIT distance="650" swimtime="00:09:17.26" />
                    <SPLIT distance="700" swimtime="00:10:00.60" />
                    <SPLIT distance="750" swimtime="00:10:42.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="390" swimtime="00:01:27.76" resultid="8074" heatid="10586" lane="2" entrytime="00:01:28.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="332" swimtime="00:02:41.99" resultid="8075" heatid="10656" lane="1" entrytime="00:02:35.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.05" />
                    <SPLIT distance="100" swimtime="00:01:17.87" />
                    <SPLIT distance="150" swimtime="00:02:00.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Steven" lastname="Matheussi Viana E Silva" birthdate="2012-05-03" gender="M" nation="BRA" license="376986" swrid="5588810" athleteid="8284" externalid="376986">
              <RESULTS>
                <RESULT eventid="1087" points="366" swimtime="00:02:55.37" resultid="8285" heatid="10490" lane="1" entrytime="00:02:56.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                    <SPLIT distance="100" swimtime="00:01:23.63" />
                    <SPLIT distance="150" swimtime="00:02:08.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="352" swimtime="00:01:05.66" resultid="8286" heatid="10541" lane="5" entrytime="00:01:10.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="342" swimtime="00:01:21.31" resultid="8287" heatid="10596" lane="9" entrytime="00:01:20.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="321" swimtime="00:02:46.38" resultid="8288" heatid="10648" lane="2" entrytime="00:02:51.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.69" />
                    <SPLIT distance="100" swimtime="00:01:23.03" />
                    <SPLIT distance="150" swimtime="00:02:08.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="252" swimtime="00:01:18.28" resultid="8289" heatid="10706" lane="9" entrytime="00:01:20.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinícius" lastname="Oliveira Cruz" birthdate="2005-07-02" gender="M" nation="BRA" license="298495" swrid="5653299" athleteid="8351" externalid="298495" level="ADTRISC">
              <RESULTS>
                <RESULT eventid="1289" points="740" swimtime="00:01:52.76" resultid="8352" heatid="10674" lane="4" entrytime="00:01:50.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.62" />
                    <SPLIT distance="100" swimtime="00:00:54.59" />
                    <SPLIT distance="150" swimtime="00:01:23.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olavo" lastname="Valduga Artigas" birthdate="2012-06-26" gender="M" nation="BRA" license="369270" swrid="5588941" athleteid="8169" externalid="369270">
              <RESULTS>
                <RESULT eventid="1087" points="208" swimtime="00:03:31.66" resultid="8170" heatid="10487" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.25" />
                    <SPLIT distance="100" swimtime="00:01:43.14" />
                    <SPLIT distance="150" swimtime="00:02:39.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="222" swimtime="00:01:16.58" resultid="8171" heatid="10538" lane="5" entrytime="00:01:21.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="212" swimtime="00:00:35.03" resultid="8172" heatid="10614" lane="0" entrytime="00:00:35.57" entrycourse="LCM" />
                <RESULT eventid="1219" points="174" swimtime="00:01:41.76" resultid="8173" heatid="10592" lane="8" entrytime="00:01:43.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="214" swimtime="00:03:10.31" resultid="8174" heatid="10646" lane="4" entrytime="00:03:09.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.49" />
                    <SPLIT distance="100" swimtime="00:01:39.65" />
                    <SPLIT distance="150" swimtime="00:02:32.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="240" swimtime="00:05:53.96" resultid="8175" heatid="10719" lane="8" entrytime="00:05:47.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.75" />
                    <SPLIT distance="100" swimtime="00:01:23.75" />
                    <SPLIT distance="150" swimtime="00:02:10.18" />
                    <SPLIT distance="200" swimtime="00:02:54.97" />
                    <SPLIT distance="250" swimtime="00:03:41.36" />
                    <SPLIT distance="300" swimtime="00:04:26.72" />
                    <SPLIT distance="350" swimtime="00:05:12.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Kremer De Aguiar" birthdate="2009-12-22" gender="F" nation="BRA" license="338987" swrid="5600196" athleteid="7939" externalid="338987">
              <RESULTS>
                <RESULT eventid="1079" points="420" swimtime="00:03:03.58" resultid="7940" heatid="10485" lane="8" entrytime="00:03:02.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.82" />
                    <SPLIT distance="100" swimtime="00:01:27.33" />
                    <SPLIT distance="150" swimtime="00:02:15.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="466" swimtime="00:00:37.61" resultid="7941" heatid="10565" lane="0" entrytime="00:00:37.18" entrycourse="LCM" />
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 9:12)" eventid="1211" status="DSQ" swimtime="00:01:24.39" resultid="7942" heatid="10588" lane="8" entrytime="00:01:23.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="448" swimtime="00:02:44.76" resultid="7943" heatid="10643" lane="2" entrytime="00:02:44.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                    <SPLIT distance="100" swimtime="00:01:20.24" />
                    <SPLIT distance="150" swimtime="00:02:05.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Ferreira Motta" birthdate="2008-10-24" gender="M" nation="BRA" license="378068" swrid="5600160" athleteid="8290" externalid="378068">
              <RESULTS>
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="8291" heatid="10574" lane="1" entrytime="00:00:34.54" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabio" lastname="Chiquito Do Brasil" birthdate="2011-05-11" gender="M" nation="BRA" license="413921" swrid="5811240" athleteid="8366" externalid="413921">
              <RESULTS>
                <RESULT eventid="1123" points="357" swimtime="00:10:37.24" resultid="8367" heatid="10517" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                    <SPLIT distance="100" swimtime="00:01:14.53" />
                    <SPLIT distance="150" swimtime="00:01:54.38" />
                    <SPLIT distance="200" swimtime="00:02:34.59" />
                    <SPLIT distance="250" swimtime="00:03:14.90" />
                    <SPLIT distance="300" swimtime="00:03:55.25" />
                    <SPLIT distance="350" swimtime="00:04:35.78" />
                    <SPLIT distance="400" swimtime="00:05:16.21" />
                    <SPLIT distance="450" swimtime="00:05:56.60" />
                    <SPLIT distance="500" swimtime="00:06:37.22" />
                    <SPLIT distance="550" swimtime="00:07:17.65" />
                    <SPLIT distance="600" swimtime="00:07:58.29" />
                    <SPLIT distance="650" swimtime="00:08:38.51" />
                    <SPLIT distance="700" swimtime="00:09:18.94" />
                    <SPLIT distance="750" swimtime="00:09:58.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="380" swimtime="00:01:04.01" resultid="8368" heatid="10535" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="386" swimtime="00:00:28.69" resultid="8369" heatid="10619" lane="2" entrytime="00:00:29.87" entrycourse="LCM" />
                <RESULT eventid="1289" points="415" swimtime="00:02:16.65" resultid="8370" heatid="10663" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.55" />
                    <SPLIT distance="100" swimtime="00:01:06.27" />
                    <SPLIT distance="150" swimtime="00:01:41.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="405" swimtime="00:04:57.31" resultid="8371" heatid="10720" lane="6" entrytime="00:05:03.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                    <SPLIT distance="100" swimtime="00:01:08.86" />
                    <SPLIT distance="150" swimtime="00:01:45.80" />
                    <SPLIT distance="200" swimtime="00:02:23.43" />
                    <SPLIT distance="250" swimtime="00:03:01.96" />
                    <SPLIT distance="300" swimtime="00:03:41.00" />
                    <SPLIT distance="350" swimtime="00:04:20.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="295" swimtime="00:01:17.47" resultid="8372" heatid="10735" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorena" lastname="Mascarenhas" birthdate="2011-08-31" gender="F" nation="BRA" license="370581" swrid="5602558" athleteid="8242" externalid="370581">
              <RESULTS>
                <RESULT eventid="1063" points="433" swimtime="00:02:42.71" resultid="8243" heatid="10472" lane="5" entrytime="00:02:45.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                    <SPLIT distance="100" swimtime="00:01:18.70" />
                    <SPLIT distance="150" swimtime="00:02:01.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="452" swimtime="00:01:07.36" resultid="8244" heatid="10530" lane="5" entrytime="00:01:08.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="408" swimtime="00:00:31.81" resultid="8245" heatid="10604" lane="5" entrytime="00:00:31.90" entrycourse="LCM" />
                <RESULT eventid="1211" points="359" swimtime="00:01:30.21" resultid="8246" heatid="10586" lane="9" entrytime="00:01:31.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="414" swimtime="00:02:49.12" resultid="8247" heatid="10642" lane="3" entrytime="00:02:49.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                    <SPLIT distance="100" swimtime="00:01:21.67" />
                    <SPLIT distance="150" swimtime="00:02:11.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="440" swimtime="00:01:15.08" resultid="8248" heatid="10732" lane="9" entrytime="00:01:14.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Kirchgassner" birthdate="2007-02-10" gender="M" nation="BRA" license="313535" swrid="5600230" athleteid="7898" externalid="313535">
              <RESULTS>
                <RESULT eventid="1187" points="611" swimtime="00:00:30.58" resultid="7899" heatid="10575" lane="0" entrytime="00:00:31.14" entrycourse="LCM" />
                <RESULT eventid="1219" points="670" swimtime="00:01:04.98" resultid="7900" heatid="10599" lane="3" entrytime="00:01:04.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Garcia De Fraga" birthdate="2009-03-24" gender="M" nation="BRA" license="342147" swrid="5600172" athleteid="7840" externalid="342147">
              <RESULTS>
                <RESULT eventid="1071" points="607" swimtime="00:02:12.16" resultid="7841" heatid="10480" lane="5" entrytime="00:02:12.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                    <SPLIT distance="100" swimtime="00:01:05.74" />
                    <SPLIT distance="150" swimtime="00:01:39.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="585" swimtime="00:00:55.47" resultid="7842" heatid="10551" lane="0" entrytime="00:00:56.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.29" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.5 - Pés não virados para fora durante a parte propulsora da pernada (fim do ciclo).  (Horário: 9:24)" eventid="1219" status="DSQ" swimtime="00:01:11.51" resultid="7843" heatid="10591" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="612" swimtime="00:02:14.22" resultid="7844" heatid="10652" lane="5" entrytime="00:02:15.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.22" />
                    <SPLIT distance="100" swimtime="00:01:02.30" />
                    <SPLIT distance="150" swimtime="00:01:41.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="618" swimtime="00:01:00.56" resultid="7845" heatid="10742" lane="4" entrytime="00:00:59.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Fontoura" birthdate="2010-08-26" gender="M" nation="BRA" license="338922" swrid="5600167" athleteid="8020" externalid="338922">
              <RESULTS>
                <RESULT eventid="1103" points="334" swimtime="00:00:32.07" resultid="8021" heatid="10505" lane="9" entrytime="00:00:32.60" entrycourse="LCM" />
                <RESULT eventid="1155" points="423" swimtime="00:01:01.77" resultid="8022" heatid="10546" lane="6" entrytime="00:01:02.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="398" swimtime="00:00:28.41" resultid="8023" heatid="10621" lane="1" entrytime="00:00:28.88" entrycourse="LCM" />
                <RESULT eventid="1273" points="340" swimtime="00:02:43.29" resultid="8024" heatid="10648" lane="4" entrytime="00:02:44.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:18.32" />
                    <SPLIT distance="150" swimtime="00:02:07.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="359" swimtime="00:02:23.46" resultid="8025" heatid="10668" lane="6" entrytime="00:02:21.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                    <SPLIT distance="100" swimtime="00:01:08.93" />
                    <SPLIT distance="150" swimtime="00:01:46.32" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 9:19), Na volta dos 50m." eventid="1341" status="DSQ" swimtime="00:01:12.06" resultid="8026" heatid="10707" lane="8" entrytime="00:01:14.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="16" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1205" points="606" swimtime="00:08:14.50" resultid="8419" heatid="10580" lane="2" entrytime="00:08:10.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.18" />
                    <SPLIT distance="100" swimtime="00:00:59.04" />
                    <SPLIT distance="150" swimtime="00:01:31.11" />
                    <SPLIT distance="200" swimtime="00:02:02.44" />
                    <SPLIT distance="250" swimtime="00:02:29.88" />
                    <SPLIT distance="300" swimtime="00:03:01.66" />
                    <SPLIT distance="350" swimtime="00:03:36.70" />
                    <SPLIT distance="400" swimtime="00:04:10.62" />
                    <SPLIT distance="450" swimtime="00:04:37.76" />
                    <SPLIT distance="500" swimtime="00:05:08.36" />
                    <SPLIT distance="550" swimtime="00:05:40.15" />
                    <SPLIT distance="600" swimtime="00:06:13.93" />
                    <SPLIT distance="650" swimtime="00:06:41.88" />
                    <SPLIT distance="700" swimtime="00:07:11.94" />
                    <SPLIT distance="750" swimtime="00:07:43.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7901" number="1" />
                    <RELAYPOSITION athleteid="8307" number="2" />
                    <RELAYPOSITION athleteid="7840" number="3" />
                    <RELAYPOSITION athleteid="7884" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="19" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1207" points="610" swimtime="00:08:13.49" resultid="8420" heatid="10581" lane="5" entrytime="00:07:27.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.98" />
                    <SPLIT distance="100" swimtime="00:00:58.59" />
                    <SPLIT distance="150" swimtime="00:01:30.47" />
                    <SPLIT distance="200" swimtime="00:02:02.31" />
                    <SPLIT distance="250" swimtime="00:02:29.40" />
                    <SPLIT distance="300" swimtime="00:02:59.48" />
                    <SPLIT distance="350" swimtime="00:03:31.01" />
                    <SPLIT distance="400" swimtime="00:04:01.42" />
                    <SPLIT distance="450" swimtime="00:04:31.94" />
                    <SPLIT distance="500" swimtime="00:05:06.19" />
                    <SPLIT distance="550" swimtime="00:05:41.36" />
                    <SPLIT distance="600" swimtime="00:06:15.75" />
                    <SPLIT distance="650" swimtime="00:06:42.87" />
                    <SPLIT distance="700" swimtime="00:07:12.94" />
                    <SPLIT distance="750" swimtime="00:07:43.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7898" number="1" />
                    <RELAYPOSITION athleteid="8118" number="2" />
                    <RELAYPOSITION athleteid="8378" number="3" />
                    <RELAYPOSITION athleteid="7892" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1203" points="506" swimtime="00:08:45.19" resultid="8421" heatid="10579" lane="4" entrytime="00:08:20.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                    <SPLIT distance="100" swimtime="00:01:02.91" />
                    <SPLIT distance="150" swimtime="00:01:35.56" />
                    <SPLIT distance="200" swimtime="00:02:08.08" />
                    <SPLIT distance="250" swimtime="00:02:36.95" />
                    <SPLIT distance="300" swimtime="00:03:10.15" />
                    <SPLIT distance="350" swimtime="00:03:45.86" />
                    <SPLIT distance="400" swimtime="00:04:20.22" />
                    <SPLIT distance="450" swimtime="00:04:50.86" />
                    <SPLIT distance="500" swimtime="00:05:26.13" />
                    <SPLIT distance="550" swimtime="00:06:01.91" />
                    <SPLIT distance="600" swimtime="00:06:35.66" />
                    <SPLIT distance="650" swimtime="00:07:03.97" />
                    <SPLIT distance="700" swimtime="00:07:36.90" />
                    <SPLIT distance="750" swimtime="00:08:11.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8048" number="1" />
                    <RELAYPOSITION athleteid="8384" number="2" />
                    <RELAYPOSITION athleteid="8034" number="3" />
                    <RELAYPOSITION athleteid="8235" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1331" points="564" swimtime="00:04:10.17" resultid="8422" heatid="10698" lane="4" entrytime="00:03:51.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.80" />
                    <SPLIT distance="100" swimtime="00:01:03.03" />
                    <SPLIT distance="150" swimtime="00:01:34.81" />
                    <SPLIT distance="200" swimtime="00:02:10.51" />
                    <SPLIT distance="250" swimtime="00:02:41.14" />
                    <SPLIT distance="300" swimtime="00:03:16.24" />
                    <SPLIT distance="350" swimtime="00:03:41.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7965" number="1" />
                    <RELAYPOSITION athleteid="8266" number="2" />
                    <RELAYPOSITION athleteid="8118" number="3" />
                    <RELAYPOSITION athleteid="8337" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1399" points="640" swimtime="00:03:38.41" resultid="8427" heatid="10753" lane="4" entrytime="00:03:28.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.22" />
                    <SPLIT distance="100" swimtime="00:00:53.75" />
                    <SPLIT distance="150" swimtime="00:01:19.58" />
                    <SPLIT distance="200" swimtime="00:01:47.78" />
                    <SPLIT distance="250" swimtime="00:02:14.21" />
                    <SPLIT distance="300" swimtime="00:02:43.01" />
                    <SPLIT distance="350" swimtime="00:03:09.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8337" number="1" />
                    <RELAYPOSITION athleteid="7892" number="2" />
                    <RELAYPOSITION athleteid="8118" number="3" />
                    <RELAYPOSITION athleteid="7857" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1329" points="574" swimtime="00:04:08.67" resultid="8423" heatid="10697" lane="4" entrytime="00:04:06.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                    <SPLIT distance="100" swimtime="00:01:02.16" />
                    <SPLIT distance="150" swimtime="00:01:34.23" />
                    <SPLIT distance="200" swimtime="00:02:11.66" />
                    <SPLIT distance="250" swimtime="00:02:40.00" />
                    <SPLIT distance="300" swimtime="00:03:12.15" />
                    <SPLIT distance="350" swimtime="00:03:38.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7908" number="1" />
                    <RELAYPOSITION athleteid="8373" number="2" />
                    <RELAYPOSITION athleteid="8344" number="3" />
                    <RELAYPOSITION athleteid="7840" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1397" points="596" swimtime="00:03:43.60" resultid="8428" heatid="10752" lane="4" entrytime="00:03:37.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.32" />
                    <SPLIT distance="100" swimtime="00:00:55.23" />
                    <SPLIT distance="150" swimtime="00:01:21.50" />
                    <SPLIT distance="200" swimtime="00:01:50.51" />
                    <SPLIT distance="250" swimtime="00:02:17.80" />
                    <SPLIT distance="300" swimtime="00:02:47.64" />
                    <SPLIT distance="350" swimtime="00:03:14.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7908" number="1" />
                    <RELAYPOSITION athleteid="7840" number="2" />
                    <RELAYPOSITION athleteid="8344" number="3" />
                    <RELAYPOSITION athleteid="7884" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1323" points="360" swimtime="00:04:50.51" resultid="8424" heatid="10693" lane="4" entrytime="00:04:40.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                    <SPLIT distance="100" swimtime="00:01:08.98" />
                    <SPLIT distance="150" swimtime="00:01:46.97" />
                    <SPLIT distance="200" swimtime="00:02:29.72" />
                    <SPLIT distance="250" swimtime="00:03:04.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8384" number="1" />
                    <RELAYPOSITION athleteid="8284" number="2" />
                    <RELAYPOSITION athleteid="8215" number="3" />
                    <RELAYPOSITION athleteid="8162" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1391" points="403" swimtime="00:04:14.84" resultid="8431" heatid="10748" lane="3" entrytime="00:04:07.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.32" />
                    <SPLIT distance="100" swimtime="00:01:00.31" />
                    <SPLIT distance="150" swimtime="00:01:30.71" />
                    <SPLIT distance="200" swimtime="00:02:05.56" />
                    <SPLIT distance="250" swimtime="00:02:36.57" />
                    <SPLIT distance="350" swimtime="00:03:41.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8384" number="1" />
                    <RELAYPOSITION athleteid="8162" number="2" />
                    <RELAYPOSITION athleteid="8176" number="3" />
                    <RELAYPOSITION athleteid="8122" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1327" points="423" swimtime="00:04:35.29" resultid="8425" heatid="10696" lane="4" entrytime="00:04:09.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                    <SPLIT distance="100" swimtime="00:01:07.16" />
                    <SPLIT distance="150" swimtime="00:01:45.55" />
                    <SPLIT distance="200" swimtime="00:02:30.02" />
                    <SPLIT distance="250" swimtime="00:03:03.25" />
                    <SPLIT distance="300" swimtime="00:03:39.60" />
                    <SPLIT distance="350" swimtime="00:04:05.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7999" number="1" />
                    <RELAYPOSITION athleteid="8307" number="2" />
                    <RELAYPOSITION athleteid="8027" number="3" />
                    <RELAYPOSITION athleteid="7901" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1395" points="542" swimtime="00:03:50.79" resultid="8429" heatid="10751" lane="4" entrytime="00:03:42.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.48" />
                    <SPLIT distance="100" swimtime="00:00:56.09" />
                    <SPLIT distance="150" swimtime="00:01:22.66" />
                    <SPLIT distance="200" swimtime="00:01:53.12" />
                    <SPLIT distance="250" swimtime="00:02:20.63" />
                    <SPLIT distance="300" swimtime="00:02:51.83" />
                    <SPLIT distance="350" swimtime="00:03:20.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7901" number="1" />
                    <RELAYPOSITION athleteid="8307" number="2" />
                    <RELAYPOSITION athleteid="8013" number="3" />
                    <RELAYPOSITION athleteid="7999" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1325" points="414" swimtime="00:04:37.32" resultid="8426" heatid="10695" lane="4" entrytime="00:04:37.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.97" />
                    <SPLIT distance="100" swimtime="00:01:08.53" />
                    <SPLIT distance="150" swimtime="00:01:44.50" />
                    <SPLIT distance="200" swimtime="00:02:26.82" />
                    <SPLIT distance="250" swimtime="00:03:00.04" />
                    <SPLIT distance="300" swimtime="00:03:37.62" />
                    <SPLIT distance="350" swimtime="00:04:06.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8235" number="1" />
                    <RELAYPOSITION athleteid="8090" number="2" />
                    <RELAYPOSITION athleteid="8041" number="3" />
                    <RELAYPOSITION athleteid="8048" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1393" points="488" swimtime="00:03:59.01" resultid="8430" heatid="10750" lane="4" entrytime="00:03:52.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.02" />
                    <SPLIT distance="100" swimtime="00:00:58.36" />
                    <SPLIT distance="150" swimtime="00:01:27.05" />
                    <SPLIT distance="200" swimtime="00:01:58.56" />
                    <SPLIT distance="250" swimtime="00:02:27.61" />
                    <SPLIT distance="300" swimtime="00:02:59.62" />
                    <SPLIT distance="350" swimtime="00:03:28.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8235" number="1" />
                    <RELAYPOSITION athleteid="8090" number="2" />
                    <RELAYPOSITION athleteid="8034" number="3" />
                    <RELAYPOSITION athleteid="8048" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1329" points="509" swimtime="00:04:18.92" resultid="8443" heatid="10697" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                    <SPLIT distance="100" swimtime="00:01:05.26" />
                    <SPLIT distance="150" swimtime="00:01:39.20" />
                    <SPLIT distance="200" swimtime="00:02:17.94" />
                    <SPLIT distance="250" swimtime="00:02:46.46" />
                    <SPLIT distance="300" swimtime="00:03:20.00" />
                    <SPLIT distance="350" swimtime="00:03:47.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7959" number="1" />
                    <RELAYPOSITION athleteid="7944" number="2" />
                    <RELAYPOSITION athleteid="7884" number="3" />
                    <RELAYPOSITION athleteid="8393" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1397" points="494" swimtime="00:03:57.98" resultid="8447" heatid="10752" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.32" />
                    <SPLIT distance="100" swimtime="00:00:57.39" />
                    <SPLIT distance="150" swimtime="00:01:25.97" />
                    <SPLIT distance="200" swimtime="00:01:57.63" />
                    <SPLIT distance="250" swimtime="00:02:27.30" />
                    <SPLIT distance="300" swimtime="00:02:59.11" />
                    <SPLIT distance="350" swimtime="00:03:26.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8373" number="1" />
                    <RELAYPOSITION athleteid="7959" number="2" />
                    <RELAYPOSITION athleteid="7944" number="3" />
                    <RELAYPOSITION athleteid="8393" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1323" points="290" swimtime="00:05:12.37" resultid="8444" heatid="10693" lane="3" entrytime="00:05:02.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                    <SPLIT distance="100" swimtime="00:01:18.87" />
                    <SPLIT distance="150" swimtime="00:01:57.09" />
                    <SPLIT distance="200" swimtime="00:02:41.76" />
                    <SPLIT distance="250" swimtime="00:03:20.42" />
                    <SPLIT distance="300" swimtime="00:04:05.39" />
                    <SPLIT distance="350" swimtime="00:04:36.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8129" number="1" />
                    <RELAYPOSITION athleteid="8176" number="2" />
                    <RELAYPOSITION athleteid="8135" number="3" />
                    <RELAYPOSITION athleteid="8209" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1391" points="344" swimtime="00:04:28.44" resultid="8450" heatid="10748" lane="5" entrytime="00:04:26.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                    <SPLIT distance="100" swimtime="00:01:06.53" />
                    <SPLIT distance="150" swimtime="00:01:38.42" />
                    <SPLIT distance="200" swimtime="00:02:13.84" />
                    <SPLIT distance="250" swimtime="00:02:45.52" />
                    <SPLIT distance="350" swimtime="00:03:53.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8129" number="1" />
                    <RELAYPOSITION athleteid="8284" number="2" />
                    <RELAYPOSITION athleteid="8209" number="3" />
                    <RELAYPOSITION athleteid="8182" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1327" points="388" swimtime="00:04:43.40" resultid="8445" heatid="10696" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                    <SPLIT distance="100" swimtime="00:01:10.63" />
                    <SPLIT distance="150" swimtime="00:01:48.07" />
                    <SPLIT distance="200" swimtime="00:02:28.78" />
                    <SPLIT distance="250" swimtime="00:03:01.77" />
                    <SPLIT distance="300" swimtime="00:03:41.65" />
                    <SPLIT distance="350" swimtime="00:04:11.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8006" number="1" />
                    <RELAYPOSITION athleteid="8013" number="2" />
                    <RELAYPOSITION athleteid="7971" number="3" />
                    <RELAYPOSITION athleteid="7978" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1395" points="427" swimtime="00:04:09.88" resultid="8448" heatid="10751" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.40" />
                    <SPLIT distance="100" swimtime="00:01:01.34" />
                    <SPLIT distance="150" swimtime="00:01:31.34" />
                    <SPLIT distance="200" swimtime="00:02:02.79" />
                    <SPLIT distance="250" swimtime="00:02:34.07" />
                    <SPLIT distance="300" swimtime="00:03:08.04" />
                    <SPLIT distance="350" swimtime="00:03:37.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8027" number="1" />
                    <RELAYPOSITION athleteid="8006" number="2" />
                    <RELAYPOSITION athleteid="7978" number="3" />
                    <RELAYPOSITION athleteid="8020" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1325" points="372" swimtime="00:04:47.49" resultid="8446" heatid="10695" lane="5" entrytime="00:04:46.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                    <SPLIT distance="100" swimtime="00:01:14.02" />
                    <SPLIT distance="150" swimtime="00:01:52.40" />
                    <SPLIT distance="200" swimtime="00:02:34.32" />
                    <SPLIT distance="250" swimtime="00:03:07.66" />
                    <SPLIT distance="300" swimtime="00:03:45.42" />
                    <SPLIT distance="350" swimtime="00:04:15.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8097" number="1" />
                    <RELAYPOSITION athleteid="8277" number="2" />
                    <RELAYPOSITION athleteid="8111" number="3" />
                    <RELAYPOSITION athleteid="8034" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1393" points="400" swimtime="00:04:15.32" resultid="8449" heatid="10750" lane="5" entrytime="00:04:04.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                    <SPLIT distance="150" swimtime="00:01:33.57" />
                    <SPLIT distance="200" swimtime="00:02:06.30" />
                    <SPLIT distance="250" swimtime="00:02:38.07" />
                    <SPLIT distance="300" swimtime="00:03:12.59" />
                    <SPLIT distance="350" swimtime="00:03:42.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8366" number="1" />
                    <RELAYPOSITION athleteid="8041" number="2" />
                    <RELAYPOSITION athleteid="8292" number="3" />
                    <RELAYPOSITION athleteid="8111" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1197" points="586" swimtime="00:09:06.71" resultid="8409" heatid="10577" lane="6" entrytime="00:09:02.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.31" />
                    <SPLIT distance="100" swimtime="00:01:04.44" />
                    <SPLIT distance="150" swimtime="00:01:38.41" />
                    <SPLIT distance="200" swimtime="00:02:12.32" />
                    <SPLIT distance="250" swimtime="00:02:43.16" />
                    <SPLIT distance="300" swimtime="00:03:18.70" />
                    <SPLIT distance="350" swimtime="00:03:54.48" />
                    <SPLIT distance="400" swimtime="00:04:30.30" />
                    <SPLIT distance="450" swimtime="00:05:02.13" />
                    <SPLIT distance="500" swimtime="00:05:37.48" />
                    <SPLIT distance="550" swimtime="00:06:13.56" />
                    <SPLIT distance="600" swimtime="00:06:49.34" />
                    <SPLIT distance="650" swimtime="00:07:20.25" />
                    <SPLIT distance="700" swimtime="00:07:54.81" />
                    <SPLIT distance="750" swimtime="00:08:30.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7859" number="1" />
                    <RELAYPOSITION athleteid="7826" number="2" />
                    <RELAYPOSITION athleteid="7821" number="3" />
                    <RELAYPOSITION athleteid="7865" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1195" points="518" swimtime="00:09:29.55" resultid="8410" heatid="10576" lane="2" entrytime="00:09:26.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                    <SPLIT distance="100" swimtime="00:01:06.32" />
                    <SPLIT distance="150" swimtime="00:01:42.13" />
                    <SPLIT distance="200" swimtime="00:02:18.29" />
                    <SPLIT distance="250" swimtime="00:02:51.60" />
                    <SPLIT distance="300" swimtime="00:03:29.38" />
                    <SPLIT distance="350" swimtime="00:04:07.13" />
                    <SPLIT distance="400" swimtime="00:04:44.21" />
                    <SPLIT distance="450" swimtime="00:05:15.97" />
                    <SPLIT distance="600" swimtime="00:07:05.59" />
                    <SPLIT distance="650" swimtime="00:07:36.99" />
                    <SPLIT distance="700" swimtime="00:08:14.64" />
                    <SPLIT distance="750" swimtime="00:08:53.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8149" number="1" />
                    <RELAYPOSITION athleteid="8104" number="2" />
                    <RELAYPOSITION athleteid="8142" number="3" />
                    <RELAYPOSITION athleteid="8062" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1315" points="427" swimtime="00:05:04.74" resultid="8411" heatid="10689" lane="6" entrytime="00:04:58.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.69" />
                    <SPLIT distance="100" swimtime="00:01:15.47" />
                    <SPLIT distance="150" swimtime="00:01:53.97" />
                    <SPLIT distance="200" swimtime="00:02:35.95" />
                    <SPLIT distance="250" swimtime="00:03:13.29" />
                    <SPLIT distance="300" swimtime="00:03:58.84" />
                    <SPLIT distance="350" swimtime="00:04:29.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8242" number="1" />
                    <RELAYPOSITION athleteid="8062" number="2" />
                    <RELAYPOSITION athleteid="8083" number="3" />
                    <RELAYPOSITION athleteid="8076" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1383" points="483" swimtime="00:04:24.96" resultid="8418" heatid="10744" lane="4" entrytime="00:04:22.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                    <SPLIT distance="100" swimtime="00:01:06.49" />
                    <SPLIT distance="150" swimtime="00:01:37.83" />
                    <SPLIT distance="200" swimtime="00:02:12.40" />
                    <SPLIT distance="250" swimtime="00:02:43.92" />
                    <SPLIT distance="300" swimtime="00:03:18.70" />
                    <SPLIT distance="350" swimtime="00:03:49.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8104" number="1" />
                    <RELAYPOSITION athleteid="8083" number="2" />
                    <RELAYPOSITION athleteid="8062" number="3" />
                    <RELAYPOSITION athleteid="8076" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1317" points="415" swimtime="00:05:07.74" resultid="8412" heatid="10690" lane="1" entrytime="00:04:52.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.73" />
                    <SPLIT distance="100" swimtime="00:01:17.70" />
                    <SPLIT distance="150" swimtime="00:01:56.45" />
                    <SPLIT distance="200" swimtime="00:02:40.64" />
                    <SPLIT distance="250" swimtime="00:03:18.91" />
                    <SPLIT distance="300" swimtime="00:04:04.90" />
                    <SPLIT distance="350" swimtime="00:04:34.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7985" number="1" />
                    <RELAYPOSITION athleteid="8298" number="2" />
                    <RELAYPOSITION athleteid="7871" number="3" />
                    <RELAYPOSITION athleteid="7922" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1385" points="479" swimtime="00:04:25.70" resultid="8417" heatid="10745" lane="1" entrytime="00:04:12.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.15" />
                    <SPLIT distance="100" swimtime="00:01:04.55" />
                    <SPLIT distance="150" swimtime="00:01:35.47" />
                    <SPLIT distance="200" swimtime="00:02:09.84" />
                    <SPLIT distance="250" swimtime="00:02:41.01" />
                    <SPLIT distance="300" swimtime="00:03:16.15" />
                    <SPLIT distance="350" swimtime="00:03:49.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7922" number="1" />
                    <RELAYPOSITION athleteid="7871" number="2" />
                    <RELAYPOSITION athleteid="7985" number="3" />
                    <RELAYPOSITION athleteid="7992" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1313" points="474" swimtime="00:04:54.35" resultid="8413" heatid="10688" lane="1" entrytime="00:04:52.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.27" />
                    <SPLIT distance="150" swimtime="00:01:56.82" />
                    <SPLIT distance="250" swimtime="00:03:12.22" />
                    <SPLIT distance="300" swimtime="00:03:50.63" />
                    <SPLIT distance="350" swimtime="00:04:20.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8314" number="1" />
                    <RELAYPOSITION athleteid="8189" number="2" />
                    <RELAYPOSITION athleteid="8270" number="3" />
                    <RELAYPOSITION athleteid="8149" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" points="522" swimtime="00:04:18.13" resultid="8415" heatid="10743" lane="4" entrytime="00:04:20.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                    <SPLIT distance="100" swimtime="00:01:04.79" />
                    <SPLIT distance="150" swimtime="00:01:35.46" />
                    <SPLIT distance="200" swimtime="00:02:09.07" />
                    <SPLIT distance="250" swimtime="00:02:40.05" />
                    <SPLIT distance="300" swimtime="00:03:14.56" />
                    <SPLIT distance="350" swimtime="00:03:43.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8270" number="1" />
                    <RELAYPOSITION athleteid="8142" number="2" />
                    <RELAYPOSITION athleteid="8260" number="3" />
                    <RELAYPOSITION athleteid="8149" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1319" points="520" swimtime="00:04:45.50" resultid="8414" heatid="10691" lane="4" entrytime="00:04:42.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                    <SPLIT distance="100" swimtime="00:01:12.24" />
                    <SPLIT distance="150" swimtime="00:01:49.24" />
                    <SPLIT distance="200" swimtime="00:02:31.74" />
                    <SPLIT distance="250" swimtime="00:03:03.92" />
                    <SPLIT distance="300" swimtime="00:03:41.10" />
                    <SPLIT distance="350" swimtime="00:04:10.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7865" number="1" />
                    <RELAYPOSITION athleteid="7934" number="2" />
                    <RELAYPOSITION athleteid="7859" number="3" />
                    <RELAYPOSITION athleteid="7826" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1387" points="569" swimtime="00:04:10.83" resultid="8416" heatid="10746" lane="4" entrytime="00:04:15.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                    <SPLIT distance="100" swimtime="00:01:01.75" />
                    <SPLIT distance="150" swimtime="00:01:31.13" />
                    <SPLIT distance="200" swimtime="00:02:05.85" />
                    <SPLIT distance="250" swimtime="00:02:34.78" />
                    <SPLIT distance="300" swimtime="00:03:07.27" />
                    <SPLIT distance="350" swimtime="00:03:37.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7865" number="1" />
                    <RELAYPOSITION athleteid="7826" number="2" />
                    <RELAYPOSITION athleteid="7859" number="3" />
                    <RELAYPOSITION athleteid="7949" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1315" points="388" swimtime="00:05:14.83" resultid="8437" heatid="10689" lane="8" entrytime="00:05:16.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                    <SPLIT distance="100" swimtime="00:01:16.04" />
                    <SPLIT distance="150" swimtime="00:01:57.01" />
                    <SPLIT distance="200" swimtime="00:02:43.63" />
                    <SPLIT distance="250" swimtime="00:03:23.50" />
                    <SPLIT distance="300" swimtime="00:04:07.23" />
                    <SPLIT distance="350" swimtime="00:04:39.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8323" number="1" />
                    <RELAYPOSITION athleteid="8069" number="2" />
                    <RELAYPOSITION athleteid="8104" number="3" />
                    <RELAYPOSITION athleteid="8330" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1383" points="432" swimtime="00:04:35.02" resultid="8442" heatid="10744" lane="3" entrytime="00:04:32.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                    <SPLIT distance="100" swimtime="00:01:07.14" />
                    <SPLIT distance="150" swimtime="00:01:39.53" />
                    <SPLIT distance="200" swimtime="00:02:15.65" />
                    <SPLIT distance="250" swimtime="00:02:48.05" />
                    <SPLIT distance="300" swimtime="00:03:24.06" />
                    <SPLIT distance="350" swimtime="00:03:58.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8242" number="1" />
                    <RELAYPOSITION athleteid="8323" number="2" />
                    <RELAYPOSITION athleteid="8330" number="3" />
                    <RELAYPOSITION athleteid="8069" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1313" points="417" swimtime="00:05:07.33" resultid="8438" heatid="10688" lane="2" entrytime="00:05:20.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                    <SPLIT distance="100" swimtime="00:01:17.51" />
                    <SPLIT distance="150" swimtime="00:01:56.84" />
                    <SPLIT distance="200" swimtime="00:02:43.47" />
                    <SPLIT distance="250" swimtime="00:03:19.36" />
                    <SPLIT distance="300" swimtime="00:04:01.74" />
                    <SPLIT distance="350" swimtime="00:04:32.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8260" number="1" />
                    <RELAYPOSITION athleteid="8353" number="2" />
                    <RELAYPOSITION athleteid="8202" number="3" />
                    <RELAYPOSITION athleteid="8142" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" points="455" swimtime="00:04:30.21" resultid="8440" heatid="10743" lane="5" entrytime="00:04:35.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                    <SPLIT distance="100" swimtime="00:01:05.97" />
                    <SPLIT distance="150" swimtime="00:01:37.11" />
                    <SPLIT distance="200" swimtime="00:02:12.24" />
                    <SPLIT distance="250" swimtime="00:02:45.39" />
                    <SPLIT distance="300" swimtime="00:03:23.15" />
                    <SPLIT distance="350" swimtime="00:03:55.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8353" number="1" />
                    <RELAYPOSITION athleteid="8196" number="2" />
                    <RELAYPOSITION athleteid="8314" number="3" />
                    <RELAYPOSITION athleteid="8202" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT comment="SW 10.12 - Os pés perderam contato com a plataforma de partida antes que o colega de equipe anterior tocasse a borda.  (Horário: 19:18), Na volta dos 300m." eventid="1319" status="DSQ" swimtime="00:00:00.00" resultid="8439" heatid="10691" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7949" number="1" />
                    <RELAYPOSITION athleteid="7939" number="2" />
                    <RELAYPOSITION athleteid="7878" number="3" />
                    <RELAYPOSITION athleteid="7821" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1387" points="493" swimtime="00:04:23.14" resultid="8441" heatid="10746" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                    <SPLIT distance="100" swimtime="00:01:05.15" />
                    <SPLIT distance="150" swimtime="00:01:36.59" />
                    <SPLIT distance="200" swimtime="00:02:10.82" />
                    <SPLIT distance="250" swimtime="00:02:42.75" />
                    <SPLIT distance="300" swimtime="00:03:17.34" />
                    <SPLIT distance="350" swimtime="00:03:49.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7821" number="1" />
                    <RELAYPOSITION athleteid="7878" number="2" />
                    <RELAYPOSITION athleteid="7939" number="3" />
                    <RELAYPOSITION athleteid="7934" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1113" points="447" swimtime="00:04:44.27" resultid="8432" heatid="10510" lane="4" entrytime="00:04:42.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                    <SPLIT distance="150" swimtime="00:01:45.29" />
                    <SPLIT distance="200" swimtime="00:02:27.77" />
                    <SPLIT distance="250" swimtime="00:03:00.91" />
                    <SPLIT distance="300" swimtime="00:03:39.20" />
                    <SPLIT distance="350" swimtime="00:04:09.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8235" number="1" />
                    <RELAYPOSITION athleteid="8062" number="2" />
                    <RELAYPOSITION athleteid="8041" number="3" />
                    <RELAYPOSITION athleteid="8104" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1111" points="440" swimtime="00:04:45.79" resultid="8433" heatid="10509" lane="4" entrytime="00:04:38.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                    <SPLIT distance="100" swimtime="00:01:08.92" />
                    <SPLIT distance="150" swimtime="00:01:46.08" />
                    <SPLIT distance="200" swimtime="00:02:29.81" />
                    <SPLIT distance="250" swimtime="00:03:03.10" />
                    <SPLIT distance="300" swimtime="00:03:39.84" />
                    <SPLIT distance="350" swimtime="00:04:10.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8384" number="1" />
                    <RELAYPOSITION athleteid="8189" number="2" />
                    <RELAYPOSITION athleteid="8270" number="3" />
                    <RELAYPOSITION athleteid="8162" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1247" points="476" swimtime="00:04:38.45" resultid="8434" heatid="10631" lane="4" entrytime="00:04:22.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                    <SPLIT distance="100" swimtime="00:01:03.71" />
                    <SPLIT distance="150" swimtime="00:01:41.09" />
                    <SPLIT distance="200" swimtime="00:02:24.25" />
                    <SPLIT distance="250" swimtime="00:03:01.33" />
                    <SPLIT distance="300" swimtime="00:03:44.53" />
                    <SPLIT distance="350" swimtime="00:04:09.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7965" number="1" />
                    <RELAYPOSITION athleteid="8249" number="2" />
                    <RELAYPOSITION athleteid="7855" number="3" />
                    <RELAYPOSITION athleteid="8337" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1243" points="450" swimtime="00:04:43.53" resultid="8435" heatid="10629" lane="4" entrytime="00:04:27.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.49" />
                    <SPLIT distance="150" swimtime="00:01:47.27" />
                    <SPLIT distance="200" swimtime="00:02:30.23" />
                    <SPLIT distance="250" swimtime="00:03:03.54" />
                    <SPLIT distance="300" swimtime="00:03:38.55" />
                    <SPLIT distance="350" swimtime="00:04:08.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8307" number="1" />
                    <RELAYPOSITION athleteid="7871" number="2" />
                    <RELAYPOSITION athleteid="8006" number="3" />
                    <RELAYPOSITION athleteid="7922" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1245" points="587" swimtime="00:04:19.58" resultid="8436" heatid="10630" lane="4" entrytime="00:04:22.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.18" />
                    <SPLIT distance="100" swimtime="00:01:00.71" />
                    <SPLIT distance="150" swimtime="00:01:33.07" />
                    <SPLIT distance="200" swimtime="00:02:10.67" />
                    <SPLIT distance="250" swimtime="00:02:41.51" />
                    <SPLIT distance="300" swimtime="00:03:17.41" />
                    <SPLIT distance="350" swimtime="00:03:46.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7908" number="1" />
                    <RELAYPOSITION athleteid="8373" number="2" />
                    <RELAYPOSITION athleteid="7865" number="3" />
                    <RELAYPOSITION athleteid="7826" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1113" points="408" swimtime="00:04:53.13" resultid="8451" heatid="10510" lane="6" entrytime="00:04:53.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                    <SPLIT distance="100" swimtime="00:01:16.09" />
                    <SPLIT distance="150" swimtime="00:01:52.85" />
                    <SPLIT distance="200" swimtime="00:02:34.46" />
                    <SPLIT distance="250" swimtime="00:03:07.65" />
                    <SPLIT distance="300" swimtime="00:03:46.85" />
                    <SPLIT distance="350" swimtime="00:04:18.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8242" number="1" />
                    <RELAYPOSITION athleteid="8048" number="2" />
                    <RELAYPOSITION athleteid="8034" number="3" />
                    <RELAYPOSITION athleteid="8083" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1111" points="384" swimtime="00:04:59.10" resultid="8452" heatid="10509" lane="5" entrytime="00:04:53.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                    <SPLIT distance="100" swimtime="00:01:17.73" />
                    <SPLIT distance="150" swimtime="00:01:56.61" />
                    <SPLIT distance="200" swimtime="00:02:39.68" />
                    <SPLIT distance="250" swimtime="00:03:14.47" />
                    <SPLIT distance="300" swimtime="00:03:56.17" />
                    <SPLIT distance="350" swimtime="00:04:25.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8314" number="1" />
                    <RELAYPOSITION athleteid="8284" number="2" />
                    <RELAYPOSITION athleteid="8215" number="3" />
                    <RELAYPOSITION athleteid="8149" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1243" points="416" swimtime="00:04:51.20" resultid="8453" heatid="10629" lane="6" entrytime="00:04:37.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                    <SPLIT distance="100" swimtime="00:01:17.73" />
                    <SPLIT distance="150" swimtime="00:01:57.00" />
                    <SPLIT distance="200" swimtime="00:02:41.57" />
                    <SPLIT distance="250" swimtime="00:03:16.58" />
                    <SPLIT distance="300" swimtime="00:03:55.29" />
                    <SPLIT distance="350" swimtime="00:04:22.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7985" number="1" />
                    <RELAYPOSITION athleteid="8298" number="2" />
                    <RELAYPOSITION athleteid="8020" number="3" />
                    <RELAYPOSITION athleteid="7901" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1245" points="550" swimtime="00:04:25.28" resultid="8454" heatid="10630" lane="5" entrytime="00:04:26.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                    <SPLIT distance="100" swimtime="00:01:00.92" />
                    <SPLIT distance="150" swimtime="00:01:39.13" />
                    <SPLIT distance="200" swimtime="00:02:20.58" />
                    <SPLIT distance="250" swimtime="00:02:48.45" />
                    <SPLIT distance="300" swimtime="00:03:21.53" />
                    <SPLIT distance="350" swimtime="00:03:51.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7840" number="1" />
                    <RELAYPOSITION athleteid="7934" number="2" />
                    <RELAYPOSITION athleteid="8344" number="3" />
                    <RELAYPOSITION athleteid="7949" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="16044" nation="BRA" region="SC" clubid="8838" swrid="94001" name="Instituto Coree">
          <ATHLETES>
            <ATHLETE firstname="Bruna" lastname="Mendes Costa" birthdate="2010-05-27" gender="F" nation="BRA" license="392182" swrid="5756233" athleteid="8858" externalid="392182">
              <RESULTS>
                <RESULT eventid="1063" points="390" status="EXH" swimtime="00:02:48.49" resultid="8859" heatid="10472" lane="7" entrytime="00:02:47.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.38" />
                    <SPLIT distance="100" swimtime="00:01:22.36" />
                    <SPLIT distance="150" swimtime="00:02:06.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="447" status="EXH" swimtime="00:00:30.87" resultid="8860" heatid="10605" lane="6" entrytime="00:00:31.40" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariana" lastname="Lima Acevedo" birthdate="2012-05-12" gender="F" nation="BRA" license="378153" swrid="5627284" athleteid="8851" externalid="378153">
              <RESULTS>
                <RESULT eventid="1079" points="354" status="EXH" swimtime="00:03:14.36" resultid="8852" heatid="10483" lane="3" entrytime="00:03:12.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.10" />
                    <SPLIT distance="100" swimtime="00:01:33.94" />
                    <SPLIT distance="150" swimtime="00:02:25.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="360" status="EXH" swimtime="00:06:11.54" resultid="8853" heatid="10519" lane="7" entrytime="00:06:15.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.60" />
                    <SPLIT distance="100" swimtime="00:01:32.41" />
                    <SPLIT distance="150" swimtime="00:02:22.29" />
                    <SPLIT distance="200" swimtime="00:03:10.71" />
                    <SPLIT distance="250" swimtime="00:04:01.63" />
                    <SPLIT distance="300" swimtime="00:04:51.76" />
                    <SPLIT distance="350" swimtime="00:05:32.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="354" status="EXH" swimtime="00:01:30.59" resultid="8854" heatid="10587" lane="0" entrytime="00:01:26.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="376" status="EXH" swimtime="00:02:54.73" resultid="8855" heatid="10642" lane="7" entrytime="00:02:51.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                    <SPLIT distance="100" swimtime="00:01:26.22" />
                    <SPLIT distance="150" swimtime="00:02:17.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Torres Streit" birthdate="2012-05-22" gender="M" nation="BRA" license="408715" athleteid="8863" externalid="408715">
              <RESULTS>
                <RESULT eventid="1071" points="320" status="EXH" swimtime="00:02:43.52" resultid="8864" heatid="10476" lane="4" entrytime="00:02:45.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                    <SPLIT distance="100" swimtime="00:01:19.44" />
                    <SPLIT distance="150" swimtime="00:02:01.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentino" lastname="Thoth Da Silva" birthdate="2009-08-22" gender="M" nation="BRA" license="378150" swrid="5756256" athleteid="8845" externalid="378150">
              <RESULTS>
                <RESULT eventid="1171" points="368" status="EXH" swimtime="00:02:33.94" resultid="8846" heatid="10557" lane="4" entrytime="00:02:28.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="100" swimtime="00:01:12.86" />
                    <SPLIT distance="150" swimtime="00:01:53.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="499" status="EXH" swimtime="00:00:58.47" resultid="8847" heatid="10549" lane="4" entrytime="00:00:57.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="504" status="EXH" swimtime="00:00:26.26" resultid="8848" heatid="10626" lane="1" entrytime="00:00:25.94" entrycourse="LCM" />
                <RESULT eventid="1219" points="372" status="EXH" swimtime="00:01:19.06" resultid="8849" heatid="10596" lane="7" entrytime="00:01:19.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="465" status="EXH" swimtime="00:02:27.12" resultid="8850" heatid="10650" lane="1" entrytime="00:02:33.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.42" />
                    <SPLIT distance="100" swimtime="00:01:10.09" />
                    <SPLIT distance="150" swimtime="00:01:53.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otavio" lastname="Henrique Mühlmann Provezi" lastname.en="Henrique Muhlmann Provezi" birthdate="2012-11-14" gender="M" nation="BRA" license="378160" swrid="5684568" athleteid="8856" externalid="378160">
              <RESULTS>
                <RESULT eventid="1373" points="340" status="EXH" swimtime="00:01:13.86" resultid="8857" heatid="10738" lane="8" entrytime="00:01:15.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Luis Siewert Pretto" birthdate="2012-05-03" gender="M" nation="BRA" license="401862" swrid="5684578" athleteid="8861" externalid="401862">
              <RESULTS>
                <RESULT eventid="1219" points="302" status="EXH" swimtime="00:01:24.74" resultid="8862" heatid="10595" lane="0" entrytime="00:01:24.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Saviato" birthdate="2012-01-10" gender="M" nation="BRA" license="378149" swrid="5627371" athleteid="8843" externalid="378149">
              <RESULTS>
                <RESULT eventid="1341" points="261" status="EXH" swimtime="00:01:17.31" resultid="8844" heatid="10706" lane="5" entrytime="00:01:16.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yuri" lastname="Helmann" birthdate="2012-08-26" gender="M" nation="BRA" license="378148" swrid="5684563" athleteid="8839" externalid="378148">
              <RESULTS>
                <RESULT eventid="1123" points="242" status="EXH" swimtime="00:12:04.76" resultid="8840" heatid="10516" lane="1" entrytime="00:11:44.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.69" />
                    <SPLIT distance="100" swimtime="00:01:24.52" />
                    <SPLIT distance="150" swimtime="00:02:08.48" />
                    <SPLIT distance="200" swimtime="00:02:53.81" />
                    <SPLIT distance="250" swimtime="00:03:40.73" />
                    <SPLIT distance="300" swimtime="00:04:27.17" />
                    <SPLIT distance="350" swimtime="00:05:13.45" />
                    <SPLIT distance="400" swimtime="00:06:00.16" />
                    <SPLIT distance="450" swimtime="00:06:46.03" />
                    <SPLIT distance="500" swimtime="00:07:31.98" />
                    <SPLIT distance="550" swimtime="00:08:18.53" />
                    <SPLIT distance="600" swimtime="00:09:05.01" />
                    <SPLIT distance="650" swimtime="00:09:50.64" />
                    <SPLIT distance="700" swimtime="00:10:36.15" />
                    <SPLIT distance="750" swimtime="00:11:21.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="268" status="EXH" swimtime="00:03:14.43" resultid="8841" heatid="10488" lane="3" entrytime="00:03:25.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.30" />
                    <SPLIT distance="100" swimtime="00:01:31.86" />
                    <SPLIT distance="150" swimtime="00:02:23.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="263" status="EXH" swimtime="00:06:18.04" resultid="8842" heatid="10521" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.57" />
                    <SPLIT distance="100" swimtime="00:01:33.60" />
                    <SPLIT distance="150" swimtime="00:02:24.52" />
                    <SPLIT distance="200" swimtime="00:03:14.80" />
                    <SPLIT distance="250" swimtime="00:04:05.01" />
                    <SPLIT distance="300" swimtime="00:04:56.58" />
                    <SPLIT distance="350" swimtime="00:05:38.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="36" nation="BRA" region="PR" clubid="7558" swrid="93753" name="Associação Atlética Comercial" shortname="Comercial Cascavel">
          <ATHLETES>
            <ATHLETE firstname="Gabriel" lastname="Alves Serafini" birthdate="2008-04-15" gender="M" nation="BRA" license="351644" swrid="5596867" athleteid="7711" externalid="351644">
              <RESULTS>
                <RESULT eventid="1123" points="487" swimtime="00:09:34.64" resultid="7712" heatid="10516" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.46" />
                    <SPLIT distance="100" swimtime="00:01:01.69" />
                    <SPLIT distance="150" swimtime="00:01:35.58" />
                    <SPLIT distance="200" swimtime="00:02:10.41" />
                    <SPLIT distance="250" swimtime="00:02:47.05" />
                    <SPLIT distance="300" swimtime="00:03:23.51" />
                    <SPLIT distance="350" swimtime="00:04:00.90" />
                    <SPLIT distance="400" swimtime="00:04:37.65" />
                    <SPLIT distance="450" swimtime="00:05:15.33" />
                    <SPLIT distance="500" swimtime="00:05:52.67" />
                    <SPLIT distance="550" swimtime="00:06:29.90" />
                    <SPLIT distance="600" swimtime="00:07:07.13" />
                    <SPLIT distance="650" swimtime="00:07:44.73" />
                    <SPLIT distance="700" swimtime="00:08:22.61" />
                    <SPLIT distance="750" swimtime="00:08:59.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="507" swimtime="00:02:18.30" resultid="7713" heatid="10558" lane="6" entrytime="00:02:15.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.13" />
                    <SPLIT distance="100" swimtime="00:01:02.15" />
                    <SPLIT distance="150" swimtime="00:01:38.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="509" swimtime="00:18:10.39" resultid="7714" heatid="10638" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                    <SPLIT distance="100" swimtime="00:01:05.70" />
                    <SPLIT distance="150" swimtime="00:01:40.63" />
                    <SPLIT distance="200" swimtime="00:02:15.81" />
                    <SPLIT distance="250" swimtime="00:02:51.23" />
                    <SPLIT distance="300" swimtime="00:03:27.10" />
                    <SPLIT distance="350" swimtime="00:04:02.90" />
                    <SPLIT distance="400" swimtime="00:04:38.78" />
                    <SPLIT distance="450" swimtime="00:05:14.58" />
                    <SPLIT distance="500" swimtime="00:05:50.89" />
                    <SPLIT distance="550" swimtime="00:06:27.05" />
                    <SPLIT distance="600" swimtime="00:07:04.00" />
                    <SPLIT distance="650" swimtime="00:07:40.07" />
                    <SPLIT distance="700" swimtime="00:08:17.67" />
                    <SPLIT distance="750" swimtime="00:08:54.10" />
                    <SPLIT distance="800" swimtime="00:09:31.87" />
                    <SPLIT distance="850" swimtime="00:10:08.41" />
                    <SPLIT distance="900" swimtime="00:10:45.43" />
                    <SPLIT distance="950" swimtime="00:11:22.14" />
                    <SPLIT distance="1000" swimtime="00:11:58.89" />
                    <SPLIT distance="1050" swimtime="00:12:35.49" />
                    <SPLIT distance="1100" swimtime="00:13:12.74" />
                    <SPLIT distance="1150" swimtime="00:13:50.73" />
                    <SPLIT distance="1200" swimtime="00:14:27.92" />
                    <SPLIT distance="1250" swimtime="00:15:05.91" />
                    <SPLIT distance="1300" swimtime="00:15:43.47" />
                    <SPLIT distance="1350" swimtime="00:16:21.42" />
                    <SPLIT distance="1400" swimtime="00:16:58.50" />
                    <SPLIT distance="1450" swimtime="00:17:35.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="465" swimtime="00:02:11.65" resultid="7715" heatid="10673" lane="7" entrytime="00:02:05.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.76" />
                    <SPLIT distance="100" swimtime="00:01:00.83" />
                    <SPLIT distance="150" swimtime="00:01:36.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="514" swimtime="00:01:01.70" resultid="7716" heatid="10710" lane="4" entrytime="00:01:00.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="464" swimtime="00:04:44.23" resultid="7717" heatid="10723" lane="3" entrytime="00:04:32.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                    <SPLIT distance="100" swimtime="00:01:03.09" />
                    <SPLIT distance="150" swimtime="00:01:37.76" />
                    <SPLIT distance="200" swimtime="00:02:12.89" />
                    <SPLIT distance="250" swimtime="00:02:49.13" />
                    <SPLIT distance="300" swimtime="00:03:27.60" />
                    <SPLIT distance="350" swimtime="00:04:06.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Rinaldini" birthdate="2009-04-09" gender="M" nation="BRA" license="348289" swrid="5596932" athleteid="7585" externalid="348289">
              <RESULTS>
                <RESULT eventid="1123" points="501" swimtime="00:09:28.89" resultid="7586" heatid="10513" lane="2" entrytime="00:09:03.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.88" />
                    <SPLIT distance="100" swimtime="00:01:04.58" />
                    <SPLIT distance="150" swimtime="00:01:39.17" />
                    <SPLIT distance="200" swimtime="00:02:13.41" />
                    <SPLIT distance="250" swimtime="00:02:47.98" />
                    <SPLIT distance="300" swimtime="00:03:22.75" />
                    <SPLIT distance="350" swimtime="00:03:57.56" />
                    <SPLIT distance="400" swimtime="00:04:32.71" />
                    <SPLIT distance="450" swimtime="00:05:08.96" />
                    <SPLIT distance="500" swimtime="00:05:45.87" />
                    <SPLIT distance="550" swimtime="00:06:23.02" />
                    <SPLIT distance="600" swimtime="00:06:59.99" />
                    <SPLIT distance="650" swimtime="00:07:37.27" />
                    <SPLIT distance="700" swimtime="00:08:14.89" />
                    <SPLIT distance="750" swimtime="00:08:52.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="550" swimtime="00:02:14.61" resultid="7587" heatid="10558" lane="3" entrytime="00:02:14.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.93" />
                    <SPLIT distance="100" swimtime="00:01:04.34" />
                    <SPLIT distance="150" swimtime="00:01:39.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="504" swimtime="00:05:04.69" resultid="7588" heatid="10523" lane="3" entrytime="00:04:54.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                    <SPLIT distance="100" swimtime="00:01:05.71" />
                    <SPLIT distance="150" swimtime="00:01:47.06" />
                    <SPLIT distance="200" swimtime="00:02:27.74" />
                    <SPLIT distance="250" swimtime="00:03:12.14" />
                    <SPLIT distance="300" swimtime="00:03:57.42" />
                    <SPLIT distance="350" swimtime="00:04:31.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="505" swimtime="00:18:13.22" resultid="7589" heatid="10635" lane="2" entrytime="00:17:27.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.55" />
                    <SPLIT distance="100" swimtime="00:01:06.87" />
                    <SPLIT distance="150" swimtime="00:01:42.66" />
                    <SPLIT distance="200" swimtime="00:02:18.50" />
                    <SPLIT distance="250" swimtime="00:02:54.44" />
                    <SPLIT distance="300" swimtime="00:03:30.68" />
                    <SPLIT distance="350" swimtime="00:04:06.70" />
                    <SPLIT distance="400" swimtime="00:04:43.01" />
                    <SPLIT distance="450" swimtime="00:05:19.43" />
                    <SPLIT distance="500" swimtime="00:05:56.53" />
                    <SPLIT distance="550" swimtime="00:06:33.11" />
                    <SPLIT distance="600" swimtime="00:07:09.74" />
                    <SPLIT distance="650" swimtime="00:07:46.48" />
                    <SPLIT distance="700" swimtime="00:08:23.46" />
                    <SPLIT distance="750" swimtime="00:09:00.55" />
                    <SPLIT distance="800" swimtime="00:09:37.69" />
                    <SPLIT distance="850" swimtime="00:10:14.95" />
                    <SPLIT distance="900" swimtime="00:10:52.04" />
                    <SPLIT distance="950" swimtime="00:11:29.63" />
                    <SPLIT distance="1000" swimtime="00:12:06.95" />
                    <SPLIT distance="1050" swimtime="00:12:44.60" />
                    <SPLIT distance="1100" swimtime="00:13:22.20" />
                    <SPLIT distance="1150" swimtime="00:13:59.71" />
                    <SPLIT distance="1200" swimtime="00:14:37.59" />
                    <SPLIT distance="1250" swimtime="00:15:15.61" />
                    <SPLIT distance="1300" swimtime="00:15:52.38" />
                    <SPLIT distance="1350" swimtime="00:16:28.53" />
                    <SPLIT distance="1400" swimtime="00:17:04.13" />
                    <SPLIT distance="1450" swimtime="00:17:39.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="484" swimtime="00:02:25.13" resultid="7590" heatid="10645" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.29" />
                    <SPLIT distance="150" swimtime="00:01:52.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="557" swimtime="00:04:27.41" resultid="7591" heatid="10724" lane="1" entrytime="00:04:23.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.15" />
                    <SPLIT distance="100" swimtime="00:01:02.86" />
                    <SPLIT distance="150" swimtime="00:01:36.76" />
                    <SPLIT distance="200" swimtime="00:02:11.03" />
                    <SPLIT distance="250" swimtime="00:02:45.54" />
                    <SPLIT distance="300" swimtime="00:03:20.29" />
                    <SPLIT distance="350" swimtime="00:03:54.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Schneider Paz" birthdate="2010-04-21" gender="M" nation="BRA" license="412900" swrid="5754746" athleteid="7788" externalid="412900">
              <RESULTS>
                <RESULT eventid="1087" points="201" swimtime="00:03:33.90" resultid="7789" heatid="10487" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.48" />
                    <SPLIT distance="100" swimtime="00:01:41.09" />
                    <SPLIT distance="150" swimtime="00:02:38.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="7790" heatid="10570" lane="9" />
                <RESULT eventid="1155" points="266" swimtime="00:01:12.07" resultid="7791" heatid="10536" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="278" swimtime="00:00:32.01" resultid="7792" heatid="10611" lane="4" />
                <RESULT eventid="1219" points="191" swimtime="00:01:38.67" resultid="7793" heatid="10591" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="222" swimtime="00:02:48.22" resultid="7794" heatid="10664" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                    <SPLIT distance="100" swimtime="00:01:19.45" />
                    <SPLIT distance="150" swimtime="00:02:05.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Mariotti De Castro" birthdate="2008-06-27" gender="M" nation="BRA" license="329200" swrid="5596912" athleteid="7571" externalid="329200">
              <RESULTS>
                <RESULT eventid="1103" points="556" swimtime="00:00:27.07" resultid="7572" heatid="10502" lane="6" />
                <RESULT eventid="1071" points="533" swimtime="00:02:17.98" resultid="7573" heatid="10480" lane="1" entrytime="00:02:19.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                    <SPLIT distance="100" swimtime="00:01:07.83" />
                    <SPLIT distance="150" swimtime="00:01:43.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="583" swimtime="00:04:50.23" resultid="7574" heatid="10523" lane="4" entrytime="00:04:40.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                    <SPLIT distance="100" swimtime="00:01:02.60" />
                    <SPLIT distance="150" swimtime="00:01:40.64" />
                    <SPLIT distance="200" swimtime="00:02:18.85" />
                    <SPLIT distance="250" swimtime="00:03:02.60" />
                    <SPLIT distance="300" swimtime="00:03:44.28" />
                    <SPLIT distance="350" swimtime="00:04:17.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="510" swimtime="00:00:26.17" resultid="7575" heatid="10613" lane="7" />
                <RESULT eventid="1273" points="600" swimtime="00:02:15.09" resultid="7576" heatid="10652" lane="4" entrytime="00:02:15.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.22" />
                    <SPLIT distance="100" swimtime="00:01:04.21" />
                    <SPLIT distance="150" swimtime="00:01:45.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="586" swimtime="00:00:59.08" resultid="7577" heatid="10704" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Danilo" lastname="Rodrigues" birthdate="2011-05-23" gender="M" nation="BRA" license="370763" swrid="5596934" athleteid="7662" externalid="370763">
              <RESULTS>
                <RESULT eventid="1087" points="348" swimtime="00:02:58.29" resultid="7663" heatid="10490" lane="9" entrytime="00:02:58.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.00" />
                    <SPLIT distance="100" swimtime="00:01:25.43" />
                    <SPLIT distance="150" swimtime="00:02:12.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="347" swimtime="00:02:37.00" resultid="7664" heatid="10557" lane="2" entrytime="00:02:33.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                    <SPLIT distance="100" swimtime="00:01:15.82" />
                    <SPLIT distance="150" swimtime="00:01:56.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="389" swimtime="00:05:32.19" resultid="7665" heatid="10522" lane="1" entrytime="00:05:29.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                    <SPLIT distance="100" swimtime="00:01:14.90" />
                    <SPLIT distance="150" swimtime="00:02:00.19" />
                    <SPLIT distance="200" swimtime="00:02:44.72" />
                    <SPLIT distance="250" swimtime="00:03:30.71" />
                    <SPLIT distance="300" swimtime="00:04:18.80" />
                    <SPLIT distance="350" swimtime="00:04:56.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="372" swimtime="00:02:38.51" resultid="7666" heatid="10648" lane="3" entrytime="00:02:47.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                    <SPLIT distance="100" swimtime="00:01:16.93" />
                    <SPLIT distance="150" swimtime="00:02:03.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="348" swimtime="00:01:10.24" resultid="7667" heatid="10708" lane="7" entrytime="00:01:10.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="394" swimtime="00:05:00.15" resultid="7668" heatid="10718" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.06" />
                    <SPLIT distance="100" swimtime="00:01:10.60" />
                    <SPLIT distance="150" swimtime="00:01:49.71" />
                    <SPLIT distance="200" swimtime="00:02:28.65" />
                    <SPLIT distance="250" swimtime="00:03:07.49" />
                    <SPLIT distance="300" swimtime="00:03:46.45" />
                    <SPLIT distance="350" swimtime="00:04:24.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Cordeiro Silva" birthdate="2011-09-04" gender="M" nation="BRA" license="380664" swrid="5596877" athleteid="7683" externalid="380664">
              <RESULTS>
                <RESULT eventid="1087" points="347" swimtime="00:02:58.42" resultid="7684" heatid="10489" lane="7" entrytime="00:03:09.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.03" />
                    <SPLIT distance="100" swimtime="00:01:24.45" />
                    <SPLIT distance="150" swimtime="00:02:11.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="318" swimtime="00:00:38.01" resultid="7685" heatid="10571" lane="5" entrytime="00:00:40.96" entrycourse="LCM" />
                <RESULT eventid="1219" points="321" swimtime="00:01:23.03" resultid="7686" heatid="10594" lane="3" entrytime="00:01:26.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="305" swimtime="00:02:49.28" resultid="7687" heatid="10647" lane="7" entrytime="00:02:57.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.13" />
                    <SPLIT distance="100" swimtime="00:01:24.00" />
                    <SPLIT distance="150" swimtime="00:02:10.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="190" swimtime="00:01:25.91" resultid="7688" heatid="10703" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="225" swimtime="00:01:24.76" resultid="7689" heatid="10734" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Stein Duarte" birthdate="2010-10-03" gender="F" nation="BRA" license="351635" swrid="5588923" athleteid="7592" externalid="351635">
              <RESULTS>
                <RESULT eventid="1095" points="327" swimtime="00:00:35.46" resultid="7593" heatid="10494" lane="7" />
                <RESULT eventid="1063" points="452" swimtime="00:02:40.42" resultid="7594" heatid="10473" lane="6" entrytime="00:02:35.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                    <SPLIT distance="100" swimtime="00:01:16.67" />
                    <SPLIT distance="150" swimtime="00:01:59.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="364" swimtime="00:01:12.42" resultid="7595" heatid="10529" lane="1" entrytime="00:01:11.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="405" swimtime="00:00:31.91" resultid="7596" heatid="10601" lane="0" />
                <RESULT eventid="1297" points="459" swimtime="00:00:34.82" resultid="7597" heatid="10680" lane="7" entrytime="00:00:34.70" entrycourse="LCM" />
                <RESULT eventid="1365" points="445" swimtime="00:01:14.81" resultid="7598" heatid="10732" lane="7" entrytime="00:01:12.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Vitoria Gugel" birthdate="2011-12-08" gender="F" nation="BRA" license="365490" swrid="5588960" athleteid="7760" externalid="365490">
              <RESULTS>
                <RESULT eventid="1079" points="310" swimtime="00:03:23.10" resultid="7761" heatid="10483" lane="2" entrytime="00:03:15.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.80" />
                    <SPLIT distance="100" swimtime="00:01:38.42" />
                    <SPLIT distance="150" swimtime="00:02:32.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="251" swimtime="00:03:13.08" resultid="7762" heatid="10554" lane="8" entrytime="00:03:04.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.89" />
                    <SPLIT distance="100" swimtime="00:01:31.02" />
                    <SPLIT distance="150" swimtime="00:02:23.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="326" swimtime="00:06:23.97" resultid="7763" heatid="10519" lane="4" entrytime="00:06:05.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.39" />
                    <SPLIT distance="100" swimtime="00:01:28.49" />
                    <SPLIT distance="150" swimtime="00:02:18.29" />
                    <SPLIT distance="200" swimtime="00:03:06.53" />
                    <SPLIT distance="250" swimtime="00:04:00.26" />
                    <SPLIT distance="300" swimtime="00:04:52.64" />
                    <SPLIT distance="350" swimtime="00:05:38.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="283" swimtime="00:01:37.57" resultid="7764" heatid="10585" lane="2" entrytime="00:01:31.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="337" swimtime="00:03:01.16" resultid="7765" heatid="10641" lane="3" entrytime="00:02:59.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.07" />
                    <SPLIT distance="100" swimtime="00:01:25.05" />
                    <SPLIT distance="150" swimtime="00:02:19.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="251" swimtime="00:01:27.43" resultid="7766" heatid="10700" lane="4" entrytime="00:01:24.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Henrique Wiebbeling" birthdate="2003-08-06" gender="M" nation="BRA" license="290420" swrid="4471225" athleteid="7559" externalid="290420">
              <RESULTS>
                <RESULT eventid="1123" points="479" swimtime="00:09:37.81" resultid="7560" heatid="10517" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.36" />
                    <SPLIT distance="100" swimtime="00:01:03.92" />
                    <SPLIT distance="150" swimtime="00:01:39.16" />
                    <SPLIT distance="200" swimtime="00:02:14.78" />
                    <SPLIT distance="250" swimtime="00:02:51.19" />
                    <SPLIT distance="300" swimtime="00:03:28.08" />
                    <SPLIT distance="350" swimtime="00:04:05.06" />
                    <SPLIT distance="400" swimtime="00:04:42.16" />
                    <SPLIT distance="450" swimtime="00:05:19.58" />
                    <SPLIT distance="500" swimtime="00:05:56.81" />
                    <SPLIT distance="550" swimtime="00:06:33.73" />
                    <SPLIT distance="600" swimtime="00:07:11.08" />
                    <SPLIT distance="650" swimtime="00:07:47.89" />
                    <SPLIT distance="700" swimtime="00:08:24.69" />
                    <SPLIT distance="750" swimtime="00:09:01.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="420" swimtime="00:02:29.34" resultid="7561" heatid="10474" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                    <SPLIT distance="150" swimtime="00:01:51.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="433" swimtime="00:01:01.32" resultid="7562" heatid="10537" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" status="WDR" swimtime="00:00:00.00" resultid="7563" heatid="10638" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Zital" birthdate="1991-05-03" gender="M" nation="BRA" license="093924" swrid="5727652" athleteid="7795" externalid="093924">
              <RESULTS>
                <RESULT eventid="1305" points="477" swimtime="00:00:30.13" resultid="7796" heatid="10687" lane="7" entrytime="00:00:29.66" entrycourse="LCM" />
                <RESULT eventid="1373" points="473" swimtime="00:01:06.19" resultid="7797" heatid="10741" lane="2" entrytime="00:01:05.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Vieira Rohnelt" birthdate="2012-05-03" gender="M" nation="BRA" license="365692" swrid="5588952" athleteid="7634" externalid="365692">
              <RESULTS>
                <RESULT eventid="1071" points="248" swimtime="00:02:57.98" resultid="7635" heatid="10475" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.81" />
                    <SPLIT distance="100" swimtime="00:01:26.40" />
                    <SPLIT distance="150" swimtime="00:02:12.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="252" swimtime="00:01:13.40" resultid="7636" heatid="10537" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="257" swimtime="00:06:20.96" resultid="7637" heatid="10521" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.96" />
                    <SPLIT distance="100" swimtime="00:01:32.29" />
                    <SPLIT distance="150" swimtime="00:02:21.74" />
                    <SPLIT distance="200" swimtime="00:03:09.63" />
                    <SPLIT distance="250" swimtime="00:04:05.05" />
                    <SPLIT distance="300" swimtime="00:04:58.90" />
                    <SPLIT distance="350" swimtime="00:05:41.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="250" swimtime="00:03:00.92" resultid="7638" heatid="10647" lane="8" entrytime="00:03:03.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.89" />
                    <SPLIT distance="100" swimtime="00:01:27.91" />
                    <SPLIT distance="150" swimtime="00:02:22.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="170" swimtime="00:01:29.21" resultid="7639" heatid="10705" lane="7" entrytime="00:01:33.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="223" swimtime="00:01:25.01" resultid="7640" heatid="10736" lane="9" entrytime="00:01:26.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Gamero Prado" birthdate="2007-05-16" gender="F" nation="BRA" license="305973" swrid="5596903" athleteid="7564" externalid="305973">
              <RESULTS>
                <RESULT eventid="1095" points="340" swimtime="00:00:34.97" resultid="7565" heatid="10498" lane="9" entrytime="00:00:33.42" entrycourse="LCM" />
                <RESULT eventid="1163" points="307" swimtime="00:03:00.54" resultid="7566" heatid="10554" lane="6" entrytime="00:02:52.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                    <SPLIT distance="100" swimtime="00:01:25.09" />
                    <SPLIT distance="150" swimtime="00:02:15.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="292" swimtime="00:12:10.39" resultid="7567" heatid="10632" lane="6" entrytime="00:10:25.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.95" />
                    <SPLIT distance="100" swimtime="00:01:20.31" />
                    <SPLIT distance="150" swimtime="00:02:06.13" />
                    <SPLIT distance="200" swimtime="00:02:53.92" />
                    <SPLIT distance="250" swimtime="00:03:42.18" />
                    <SPLIT distance="300" swimtime="00:04:30.39" />
                    <SPLIT distance="350" swimtime="00:05:17.46" />
                    <SPLIT distance="400" swimtime="00:06:04.86" />
                    <SPLIT distance="450" swimtime="00:06:50.98" />
                    <SPLIT distance="500" swimtime="00:07:35.65" />
                    <SPLIT distance="550" swimtime="00:08:21.73" />
                    <SPLIT distance="600" swimtime="00:09:08.16" />
                    <SPLIT distance="650" swimtime="00:09:52.22" />
                    <SPLIT distance="700" swimtime="00:10:37.81" />
                    <SPLIT distance="750" swimtime="00:11:23.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="354" swimtime="00:02:38.52" resultid="7568" heatid="10653" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.71" />
                    <SPLIT distance="100" swimtime="00:01:16.64" />
                    <SPLIT distance="150" swimtime="00:01:58.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="359" swimtime="00:05:31.04" resultid="7569" heatid="10712" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                    <SPLIT distance="100" swimtime="00:01:15.55" />
                    <SPLIT distance="150" swimtime="00:01:57.94" />
                    <SPLIT distance="200" swimtime="00:02:40.36" />
                    <SPLIT distance="250" swimtime="00:03:23.05" />
                    <SPLIT distance="300" swimtime="00:04:06.85" />
                    <SPLIT distance="350" swimtime="00:04:50.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="333" swimtime="00:01:19.55" resultid="7570" heatid="10702" lane="9" entrytime="00:01:15.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Sehn Uren" birthdate="2009-10-15" gender="F" nation="BRA" license="357159" swrid="5596937" athleteid="7599" externalid="357159">
              <RESULTS>
                <RESULT eventid="1063" points="425" swimtime="00:02:43.72" resultid="7600" heatid="10472" lane="1" entrytime="00:02:47.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                    <SPLIT distance="100" swimtime="00:01:20.61" />
                    <SPLIT distance="150" swimtime="00:02:01.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="402" swimtime="00:05:58.03" resultid="7601" heatid="10520" lane="0" entrytime="00:06:00.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.80" />
                    <SPLIT distance="100" swimtime="00:01:29.05" />
                    <SPLIT distance="150" swimtime="00:02:14.41" />
                    <SPLIT distance="200" swimtime="00:02:58.64" />
                    <SPLIT distance="250" swimtime="00:03:48.42" />
                    <SPLIT distance="300" swimtime="00:04:36.72" />
                    <SPLIT distance="350" swimtime="00:05:18.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="401" swimtime="00:01:26.96" resultid="7602" heatid="10586" lane="7" entrytime="00:01:28.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="444" swimtime="00:02:45.25" resultid="7603" heatid="10643" lane="3" entrytime="00:02:44.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                    <SPLIT distance="100" swimtime="00:01:18.96" />
                    <SPLIT distance="150" swimtime="00:02:07.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="278" swimtime="00:01:24.49" resultid="7604" heatid="10699" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="393" swimtime="00:01:17.98" resultid="7605" heatid="10731" lane="0" entrytime="00:01:17.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emanuel" lastname="Ranieri" birthdate="2011-01-24" gender="M" nation="BRA" license="390838" swrid="5596930" athleteid="7725" externalid="390838">
              <RESULTS>
                <RESULT eventid="1071" points="362" swimtime="00:02:36.93" resultid="7726" heatid="10476" lane="6" entrytime="00:02:47.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                    <SPLIT distance="100" swimtime="00:01:15.41" />
                    <SPLIT distance="150" swimtime="00:01:56.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="387" swimtime="00:01:03.62" resultid="7727" heatid="10536" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="390" swimtime="00:05:31.75" resultid="7728" heatid="10522" lane="0" entrytime="00:05:41.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.81" />
                    <SPLIT distance="100" swimtime="00:01:16.47" />
                    <SPLIT distance="150" swimtime="00:01:59.04" />
                    <SPLIT distance="200" swimtime="00:02:40.87" />
                    <SPLIT distance="250" swimtime="00:03:29.66" />
                    <SPLIT distance="300" swimtime="00:04:19.49" />
                    <SPLIT distance="350" swimtime="00:04:56.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="383" swimtime="00:02:36.94" resultid="7729" heatid="10649" lane="2" entrytime="00:02:41.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                    <SPLIT distance="100" swimtime="00:01:13.14" />
                    <SPLIT distance="150" swimtime="00:02:01.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="385" swimtime="00:02:20.11" resultid="7730" heatid="10661" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                    <SPLIT distance="100" swimtime="00:01:06.99" />
                    <SPLIT distance="150" swimtime="00:01:45.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="319" swimtime="00:01:15.46" resultid="7731" heatid="10737" lane="3" entrytime="00:01:16.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Assakura" birthdate="2010-06-29" gender="F" nation="BRA" license="376473" swrid="5596868" athleteid="7697" externalid="376473">
              <RESULTS>
                <RESULT eventid="1079" points="527" swimtime="00:02:50.24" resultid="7698" heatid="10486" lane="8" entrytime="00:02:55.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.84" />
                    <SPLIT distance="100" swimtime="00:01:21.33" />
                    <SPLIT distance="150" swimtime="00:02:06.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="461" swimtime="00:05:42.07" resultid="7699" heatid="10520" lane="3" entrytime="00:05:45.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                    <SPLIT distance="100" swimtime="00:01:20.09" />
                    <SPLIT distance="150" swimtime="00:02:05.46" />
                    <SPLIT distance="200" swimtime="00:02:49.33" />
                    <SPLIT distance="250" swimtime="00:03:36.91" />
                    <SPLIT distance="300" swimtime="00:04:22.98" />
                    <SPLIT distance="350" swimtime="00:05:03.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="450" swimtime="00:10:32.17" resultid="7700" heatid="10634" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                    <SPLIT distance="100" swimtime="00:01:12.42" />
                    <SPLIT distance="150" swimtime="00:01:50.80" />
                    <SPLIT distance="200" swimtime="00:02:30.01" />
                    <SPLIT distance="250" swimtime="00:03:10.14" />
                    <SPLIT distance="300" swimtime="00:03:50.57" />
                    <SPLIT distance="350" swimtime="00:04:31.26" />
                    <SPLIT distance="400" swimtime="00:05:11.57" />
                    <SPLIT distance="450" swimtime="00:05:52.50" />
                    <SPLIT distance="500" swimtime="00:06:32.89" />
                    <SPLIT distance="550" swimtime="00:07:13.59" />
                    <SPLIT distance="600" swimtime="00:07:54.39" />
                    <SPLIT distance="650" swimtime="00:08:34.92" />
                    <SPLIT distance="700" swimtime="00:09:14.68" />
                    <SPLIT distance="750" swimtime="00:09:54.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="472" swimtime="00:01:22.33" resultid="7701" heatid="10588" lane="9" entrytime="00:01:23.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="480" swimtime="00:02:40.99" resultid="7702" heatid="10644" lane="1" entrytime="00:02:41.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                    <SPLIT distance="100" swimtime="00:01:17.22" />
                    <SPLIT distance="150" swimtime="00:02:02.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="466" swimtime="00:05:03.48" resultid="7703" heatid="10715" lane="1" entrytime="00:05:09.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                    <SPLIT distance="100" swimtime="00:01:10.47" />
                    <SPLIT distance="150" swimtime="00:01:49.07" />
                    <SPLIT distance="200" swimtime="00:02:28.52" />
                    <SPLIT distance="250" swimtime="00:03:07.82" />
                    <SPLIT distance="300" swimtime="00:03:47.13" />
                    <SPLIT distance="350" swimtime="00:04:25.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laisa" lastname="Bernardini" birthdate="2012-06-25" gender="F" nation="BRA" license="390843" swrid="5596872" athleteid="7732" externalid="390843">
              <RESULTS>
                <RESULT eventid="1079" points="273" swimtime="00:03:31.91" resultid="7733" heatid="10481" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.23" />
                    <SPLIT distance="100" swimtime="00:01:43.56" />
                    <SPLIT distance="150" swimtime="00:02:38.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="257" swimtime="00:00:45.86" resultid="7734" heatid="10562" lane="1" entrytime="00:00:47.42" entrycourse="LCM" />
                <RESULT eventid="1131" points="310" swimtime="00:06:30.57" resultid="7735" heatid="10518" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.84" />
                    <SPLIT distance="100" swimtime="00:01:38.49" />
                    <SPLIT distance="150" swimtime="00:02:26.83" />
                    <SPLIT distance="200" swimtime="00:03:15.68" />
                    <SPLIT distance="250" swimtime="00:04:10.09" />
                    <SPLIT distance="300" swimtime="00:05:04.36" />
                    <SPLIT distance="350" swimtime="00:05:48.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="293" swimtime="00:01:36.46" resultid="7736" heatid="10584" lane="8" entrytime="00:01:41.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="323" swimtime="00:03:03.81" resultid="7737" heatid="10640" lane="5" entrytime="00:03:11.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.26" />
                    <SPLIT distance="100" swimtime="00:01:30.65" />
                    <SPLIT distance="150" swimtime="00:02:23.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="268" swimtime="00:01:28.54" resultid="7738" heatid="10728" lane="9" entrytime="00:01:30.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Pedro Serafini" birthdate="2012-05-15" gender="M" nation="BRA" license="365488" swrid="5596924" athleteid="7718" externalid="365488">
              <RESULTS>
                <RESULT eventid="1123" points="344" swimtime="00:10:44.98" resultid="7719" heatid="10517" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:15.27" />
                    <SPLIT distance="150" swimtime="00:01:56.10" />
                    <SPLIT distance="200" swimtime="00:02:36.78" />
                    <SPLIT distance="250" swimtime="00:03:17.62" />
                    <SPLIT distance="300" swimtime="00:03:58.97" />
                    <SPLIT distance="350" swimtime="00:04:40.01" />
                    <SPLIT distance="400" swimtime="00:05:21.79" />
                    <SPLIT distance="450" swimtime="00:06:03.08" />
                    <SPLIT distance="500" swimtime="00:06:44.42" />
                    <SPLIT distance="550" swimtime="00:07:25.21" />
                    <SPLIT distance="600" swimtime="00:08:06.71" />
                    <SPLIT distance="650" swimtime="00:08:46.67" />
                    <SPLIT distance="700" swimtime="00:09:27.44" />
                    <SPLIT distance="750" swimtime="00:10:07.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="233" swimtime="00:02:59.17" resultid="7720" heatid="10555" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                    <SPLIT distance="100" swimtime="00:01:23.57" />
                    <SPLIT distance="150" swimtime="00:02:12.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="340" swimtime="00:20:47.41" resultid="7721" heatid="10637" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.31" />
                    <SPLIT distance="100" swimtime="00:01:18.38" />
                    <SPLIT distance="150" swimtime="00:01:59.81" />
                    <SPLIT distance="200" swimtime="00:02:42.30" />
                    <SPLIT distance="250" swimtime="00:03:23.80" />
                    <SPLIT distance="300" swimtime="00:04:06.32" />
                    <SPLIT distance="350" swimtime="00:04:48.59" />
                    <SPLIT distance="400" swimtime="00:05:31.04" />
                    <SPLIT distance="450" swimtime="00:06:12.82" />
                    <SPLIT distance="500" swimtime="00:06:55.23" />
                    <SPLIT distance="550" swimtime="00:07:37.68" />
                    <SPLIT distance="600" swimtime="00:08:20.11" />
                    <SPLIT distance="650" swimtime="00:09:02.34" />
                    <SPLIT distance="700" swimtime="00:09:44.56" />
                    <SPLIT distance="750" swimtime="00:10:26.70" />
                    <SPLIT distance="800" swimtime="00:11:09.02" />
                    <SPLIT distance="850" swimtime="00:11:50.81" />
                    <SPLIT distance="900" swimtime="00:12:33.17" />
                    <SPLIT distance="950" swimtime="00:13:14.54" />
                    <SPLIT distance="1000" swimtime="00:13:56.40" />
                    <SPLIT distance="1050" swimtime="00:14:37.81" />
                    <SPLIT distance="1100" swimtime="00:15:20.05" />
                    <SPLIT distance="1150" swimtime="00:16:01.16" />
                    <SPLIT distance="1200" swimtime="00:16:42.89" />
                    <SPLIT distance="1250" swimtime="00:17:24.53" />
                    <SPLIT distance="1300" swimtime="00:18:06.56" />
                    <SPLIT distance="1350" swimtime="00:18:47.52" />
                    <SPLIT distance="1400" swimtime="00:19:29.44" />
                    <SPLIT distance="1450" swimtime="00:20:09.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="315" swimtime="00:02:29.88" resultid="7722" heatid="10666" lane="1" entrytime="00:02:39.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                    <SPLIT distance="100" swimtime="00:01:12.31" />
                    <SPLIT distance="150" swimtime="00:01:52.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="229" swimtime="00:01:20.78" resultid="7723" heatid="10705" lane="2" entrytime="00:01:29.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="337" swimtime="00:05:16.14" resultid="7724" heatid="10719" lane="1" entrytime="00:05:41.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                    <SPLIT distance="100" swimtime="00:01:13.17" />
                    <SPLIT distance="150" swimtime="00:01:53.37" />
                    <SPLIT distance="200" swimtime="00:02:34.08" />
                    <SPLIT distance="250" swimtime="00:03:14.82" />
                    <SPLIT distance="300" swimtime="00:03:56.27" />
                    <SPLIT distance="350" swimtime="00:04:37.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Zimmermann" birthdate="2010-01-19" gender="M" nation="BRA" license="357160" swrid="5588977" athleteid="7606" externalid="357160">
              <RESULTS>
                <RESULT eventid="1071" points="521" swimtime="00:02:19.08" resultid="7607" heatid="10480" lane="2" entrytime="00:02:19.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                    <SPLIT distance="100" swimtime="00:01:08.51" />
                    <SPLIT distance="150" swimtime="00:01:44.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="541" swimtime="00:00:56.92" resultid="7608" heatid="10538" lane="9" entrytime="00:02:02.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="540" swimtime="00:04:57.69" resultid="7609" heatid="10523" lane="6" entrytime="00:04:56.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                    <SPLIT distance="100" swimtime="00:01:06.99" />
                    <SPLIT distance="150" swimtime="00:01:45.30" />
                    <SPLIT distance="200" swimtime="00:02:23.21" />
                    <SPLIT distance="250" swimtime="00:03:06.52" />
                    <SPLIT distance="300" swimtime="00:03:50.86" />
                    <SPLIT distance="350" swimtime="00:04:24.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="514" swimtime="00:02:22.27" resultid="7610" heatid="10652" lane="7" entrytime="00:02:21.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                    <SPLIT distance="100" swimtime="00:01:07.17" />
                    <SPLIT distance="150" swimtime="00:01:51.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="538" swimtime="00:02:05.37" resultid="7611" heatid="10673" lane="0" entrytime="00:02:06.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.18" />
                    <SPLIT distance="100" swimtime="00:00:59.94" />
                    <SPLIT distance="150" swimtime="00:01:33.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="490" swimtime="00:01:05.44" resultid="7612" heatid="10741" lane="1" entrytime="00:01:05.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raul" lastname="Bonamigo" birthdate="2010-12-01" gender="M" nation="BRA" license="344397" swrid="5588559" athleteid="7704" externalid="344397">
              <RESULTS>
                <RESULT eventid="1123" points="493" swimtime="00:09:31.94" resultid="7705" heatid="10514" lane="4" entrytime="00:09:33.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                    <SPLIT distance="100" swimtime="00:01:07.04" />
                    <SPLIT distance="150" swimtime="00:01:42.51" />
                    <SPLIT distance="200" swimtime="00:02:18.53" />
                    <SPLIT distance="250" swimtime="00:02:54.49" />
                    <SPLIT distance="300" swimtime="00:03:30.50" />
                    <SPLIT distance="350" swimtime="00:04:06.57" />
                    <SPLIT distance="400" swimtime="00:04:43.12" />
                    <SPLIT distance="450" swimtime="00:05:19.04" />
                    <SPLIT distance="500" swimtime="00:05:54.96" />
                    <SPLIT distance="550" swimtime="00:06:31.30" />
                    <SPLIT distance="600" swimtime="00:07:08.03" />
                    <SPLIT distance="650" swimtime="00:07:43.96" />
                    <SPLIT distance="700" swimtime="00:08:20.78" />
                    <SPLIT distance="750" swimtime="00:08:56.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="459" swimtime="00:02:25.05" resultid="7706" heatid="10479" lane="6" entrytime="00:02:25.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                    <SPLIT distance="100" swimtime="00:01:10.78" />
                    <SPLIT distance="150" swimtime="00:01:48.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="438" swimtime="00:05:19.26" resultid="7707" heatid="10522" lane="3" entrytime="00:05:17.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                    <SPLIT distance="100" swimtime="00:01:13.19" />
                    <SPLIT distance="150" swimtime="00:01:54.45" />
                    <SPLIT distance="200" swimtime="00:02:33.11" />
                    <SPLIT distance="250" swimtime="00:03:20.33" />
                    <SPLIT distance="300" swimtime="00:04:08.26" />
                    <SPLIT distance="350" swimtime="00:04:44.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="515" swimtime="00:18:06.04" resultid="7708" heatid="10635" lane="0" entrytime="00:18:05.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                    <SPLIT distance="100" swimtime="00:01:08.68" />
                    <SPLIT distance="150" swimtime="00:01:44.93" />
                    <SPLIT distance="200" swimtime="00:02:21.41" />
                    <SPLIT distance="250" swimtime="00:02:57.88" />
                    <SPLIT distance="300" swimtime="00:03:34.21" />
                    <SPLIT distance="350" swimtime="00:04:10.56" />
                    <SPLIT distance="400" swimtime="00:04:47.17" />
                    <SPLIT distance="450" swimtime="00:05:23.63" />
                    <SPLIT distance="500" swimtime="00:06:00.41" />
                    <SPLIT distance="550" swimtime="00:06:36.87" />
                    <SPLIT distance="600" swimtime="00:07:13.17" />
                    <SPLIT distance="650" swimtime="00:07:49.86" />
                    <SPLIT distance="700" swimtime="00:08:26.10" />
                    <SPLIT distance="750" swimtime="00:09:02.63" />
                    <SPLIT distance="800" swimtime="00:09:39.03" />
                    <SPLIT distance="850" swimtime="00:10:15.10" />
                    <SPLIT distance="900" swimtime="00:10:51.83" />
                    <SPLIT distance="950" swimtime="00:11:27.78" />
                    <SPLIT distance="1000" swimtime="00:12:04.32" />
                    <SPLIT distance="1050" swimtime="00:12:40.27" />
                    <SPLIT distance="1100" swimtime="00:13:16.29" />
                    <SPLIT distance="1150" swimtime="00:13:52.54" />
                    <SPLIT distance="1200" swimtime="00:14:29.01" />
                    <SPLIT distance="1250" swimtime="00:15:05.65" />
                    <SPLIT distance="1300" swimtime="00:15:42.36" />
                    <SPLIT distance="1350" swimtime="00:16:18.76" />
                    <SPLIT distance="1400" swimtime="00:16:55.18" />
                    <SPLIT distance="1450" swimtime="00:17:30.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="428" swimtime="00:02:31.19" resultid="7709" heatid="10651" lane="0" entrytime="00:02:29.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                    <SPLIT distance="100" swimtime="00:01:11.15" />
                    <SPLIT distance="150" swimtime="00:01:57.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="488" swimtime="00:04:39.46" resultid="7710" heatid="10722" lane="6" entrytime="00:04:43.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                    <SPLIT distance="100" swimtime="00:01:05.25" />
                    <SPLIT distance="150" swimtime="00:01:40.63" />
                    <SPLIT distance="200" swimtime="00:02:16.35" />
                    <SPLIT distance="250" swimtime="00:02:51.78" />
                    <SPLIT distance="300" swimtime="00:03:28.75" />
                    <SPLIT distance="350" swimtime="00:04:04.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Luisa Lottermann" birthdate="2011-08-26" gender="F" nation="BRA" license="382238" swrid="5596909" athleteid="7690" externalid="382238">
              <RESULTS>
                <RESULT eventid="1079" points="400" swimtime="00:03:06.62" resultid="7691" heatid="10484" lane="5" entrytime="00:03:04.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.33" />
                    <SPLIT distance="100" swimtime="00:01:30.33" />
                    <SPLIT distance="150" swimtime="00:02:18.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="257" swimtime="00:03:11.58" resultid="7692" heatid="10554" lane="0" entrytime="00:03:14.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.07" />
                    <SPLIT distance="100" swimtime="00:01:31.71" />
                    <SPLIT distance="150" swimtime="00:02:21.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="357" swimtime="00:06:12.52" resultid="7693" heatid="10519" lane="6" entrytime="00:06:10.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.79" />
                    <SPLIT distance="100" swimtime="00:01:29.54" />
                    <SPLIT distance="150" swimtime="00:02:22.72" />
                    <SPLIT distance="200" swimtime="00:03:13.54" />
                    <SPLIT distance="250" swimtime="00:04:01.48" />
                    <SPLIT distance="300" swimtime="00:04:49.16" />
                    <SPLIT distance="350" swimtime="00:05:31.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="363" swimtime="00:01:29.82" resultid="7694" heatid="10586" lane="6" entrytime="00:01:28.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="335" swimtime="00:03:01.48" resultid="7695" heatid="10641" lane="8" entrytime="00:03:02.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.83" />
                    <SPLIT distance="100" swimtime="00:01:33.68" />
                    <SPLIT distance="150" swimtime="00:02:20.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="234" swimtime="00:01:29.50" resultid="7696" heatid="10700" lane="2" entrytime="00:01:29.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jordana" lastname="Rinaldini" birthdate="2004-09-13" gender="F" nation="BRA" license="342426" swrid="5596933" athleteid="7578" externalid="342426">
              <RESULTS>
                <RESULT eventid="1095" points="369" swimtime="00:00:34.04" resultid="7579" heatid="10494" lane="6" />
                <RESULT eventid="1079" points="387" swimtime="00:03:08.75" resultid="7580" heatid="10484" lane="1" entrytime="00:03:07.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                    <SPLIT distance="100" swimtime="00:01:28.14" />
                    <SPLIT distance="150" swimtime="00:02:18.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="422" swimtime="00:00:38.86" resultid="7581" heatid="10564" lane="8" entrytime="00:00:38.96" entrycourse="LCM" />
                <RESULT eventid="1211" points="401" swimtime="00:01:26.94" resultid="7582" heatid="10587" lane="2" entrytime="00:01:25.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="416" swimtime="00:02:48.90" resultid="7583" heatid="10639" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                    <SPLIT distance="100" swimtime="00:01:18.38" />
                    <SPLIT distance="150" swimtime="00:02:07.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="347" swimtime="00:01:21.29" resultid="7584" heatid="10729" lane="4" entrytime="00:01:20.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juan" lastname="Balduíno" birthdate="2009-06-24" gender="M" nation="BRA" license="370764" swrid="5596870" athleteid="7669" externalid="370764">
              <RESULTS>
                <RESULT eventid="1103" points="537" swimtime="00:00:27.39" resultid="7670" heatid="10500" lane="4" />
                <RESULT eventid="1071" points="467" swimtime="00:02:24.24" resultid="7671" heatid="10479" lane="5" entrytime="00:02:25.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                    <SPLIT distance="100" swimtime="00:01:09.85" />
                    <SPLIT distance="150" swimtime="00:01:47.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="483" swimtime="00:02:20.59" resultid="7672" heatid="10558" lane="7" entrytime="00:02:21.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.06" />
                    <SPLIT distance="100" swimtime="00:01:03.92" />
                    <SPLIT distance="150" swimtime="00:01:40.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="507" swimtime="00:05:04.05" resultid="7673" heatid="10523" lane="0" entrytime="00:05:07.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                    <SPLIT distance="100" swimtime="00:01:04.68" />
                    <SPLIT distance="150" swimtime="00:01:44.53" />
                    <SPLIT distance="200" swimtime="00:02:23.39" />
                    <SPLIT distance="250" swimtime="00:03:08.65" />
                    <SPLIT distance="300" swimtime="00:03:54.53" />
                    <SPLIT distance="350" swimtime="00:04:30.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="531" swimtime="00:02:20.74" resultid="7674" heatid="10651" lane="3" entrytime="00:02:24.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.99" />
                    <SPLIT distance="100" swimtime="00:01:05.67" />
                    <SPLIT distance="150" swimtime="00:01:48.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="519" swimtime="00:01:01.50" resultid="7675" heatid="10710" lane="5" entrytime="00:01:01.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Colaco Da Conceicao" birthdate="2011-05-25" gender="F" nation="BRA" license="369535" swrid="5588601" athleteid="7655" externalid="369535">
              <RESULTS>
                <RESULT eventid="1115" points="402" swimtime="00:20:47.15" resultid="7656" heatid="10511" lane="1" entrytime="00:20:00.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                    <SPLIT distance="100" swimtime="00:01:15.26" />
                    <SPLIT distance="150" swimtime="00:01:55.61" />
                    <SPLIT distance="200" swimtime="00:02:36.50" />
                    <SPLIT distance="250" swimtime="00:03:17.24" />
                    <SPLIT distance="300" swimtime="00:03:59.07" />
                    <SPLIT distance="350" swimtime="00:04:40.02" />
                    <SPLIT distance="400" swimtime="00:05:22.30" />
                    <SPLIT distance="450" swimtime="00:06:04.38" />
                    <SPLIT distance="500" swimtime="00:06:46.70" />
                    <SPLIT distance="550" swimtime="00:07:28.94" />
                    <SPLIT distance="600" swimtime="00:08:10.55" />
                    <SPLIT distance="650" swimtime="00:08:53.22" />
                    <SPLIT distance="700" swimtime="00:09:36.31" />
                    <SPLIT distance="750" swimtime="00:10:18.70" />
                    <SPLIT distance="800" swimtime="00:11:01.30" />
                    <SPLIT distance="850" swimtime="00:11:43.67" />
                    <SPLIT distance="900" swimtime="00:12:26.68" />
                    <SPLIT distance="950" swimtime="00:13:09.38" />
                    <SPLIT distance="1000" swimtime="00:13:51.83" />
                    <SPLIT distance="1050" swimtime="00:14:34.26" />
                    <SPLIT distance="1100" swimtime="00:15:16.18" />
                    <SPLIT distance="1150" swimtime="00:15:58.80" />
                    <SPLIT distance="1200" swimtime="00:16:41.41" />
                    <SPLIT distance="1250" swimtime="00:17:23.50" />
                    <SPLIT distance="1300" swimtime="00:18:04.96" />
                    <SPLIT distance="1350" swimtime="00:18:45.27" />
                    <SPLIT distance="1400" swimtime="00:19:27.34" />
                    <SPLIT distance="1450" swimtime="00:20:07.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="350" swimtime="00:02:54.57" resultid="7657" heatid="10469" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="410" swimtime="00:01:09.60" resultid="7658" heatid="10524" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="431" swimtime="00:10:41.37" resultid="7659" heatid="10632" lane="3" entrytime="00:10:24.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                    <SPLIT distance="100" swimtime="00:01:12.21" />
                    <SPLIT distance="150" swimtime="00:01:51.83" />
                    <SPLIT distance="200" swimtime="00:02:30.73" />
                    <SPLIT distance="250" swimtime="00:03:11.45" />
                    <SPLIT distance="300" swimtime="00:03:52.28" />
                    <SPLIT distance="350" swimtime="00:04:32.44" />
                    <SPLIT distance="400" swimtime="00:05:13.61" />
                    <SPLIT distance="450" swimtime="00:05:55.02" />
                    <SPLIT distance="500" swimtime="00:06:36.81" />
                    <SPLIT distance="550" swimtime="00:07:18.77" />
                    <SPLIT distance="600" swimtime="00:07:59.53" />
                    <SPLIT distance="650" swimtime="00:08:41.08" />
                    <SPLIT distance="700" swimtime="00:09:22.28" />
                    <SPLIT distance="750" swimtime="00:10:02.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="455" swimtime="00:02:25.89" resultid="7660" heatid="10657" lane="9" entrytime="00:02:30.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                    <SPLIT distance="100" swimtime="00:01:10.36" />
                    <SPLIT distance="150" swimtime="00:01:48.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="420" swimtime="00:05:14.11" resultid="7661" heatid="10715" lane="2" entrytime="00:05:06.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                    <SPLIT distance="100" swimtime="00:01:12.72" />
                    <SPLIT distance="150" swimtime="00:01:52.94" />
                    <SPLIT distance="200" swimtime="00:02:33.24" />
                    <SPLIT distance="250" swimtime="00:03:13.79" />
                    <SPLIT distance="300" swimtime="00:03:54.07" />
                    <SPLIT distance="350" swimtime="00:04:35.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Schneider Paz" birthdate="2011-07-03" gender="M" nation="BRA" license="412899" swrid="5754792" athleteid="7781" externalid="412899">
              <RESULTS>
                <RESULT eventid="1087" points="200" swimtime="00:03:34.40" resultid="7782" heatid="10488" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.55" />
                    <SPLIT distance="100" swimtime="00:01:44.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="218" swimtime="00:00:43.09" resultid="7783" heatid="10568" lane="4" />
                <RESULT eventid="1155" points="271" swimtime="00:01:11.67" resultid="7784" heatid="10536" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="268" swimtime="00:00:32.43" resultid="7785" heatid="10612" lane="5" />
                <RESULT eventid="1219" points="229" swimtime="00:01:32.84" resultid="7786" heatid="10591" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="253" swimtime="00:02:41.07" resultid="7787" heatid="10661" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                    <SPLIT distance="100" swimtime="00:01:13.58" />
                    <SPLIT distance="150" swimtime="00:01:56.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amanda" lastname="Borille Busetti" birthdate="2010-02-17" gender="F" nation="BRA" license="392830" swrid="5622263" athleteid="7767" externalid="392830">
              <RESULTS>
                <RESULT eventid="1063" points="304" swimtime="00:03:03.09" resultid="7768" heatid="10470" lane="2" entrytime="00:03:03.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="296" swimtime="00:06:36.62" resultid="7769" heatid="10518" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.17" />
                    <SPLIT distance="100" swimtime="00:01:34.83" />
                    <SPLIT distance="150" swimtime="00:02:28.59" />
                    <SPLIT distance="200" swimtime="00:03:20.32" />
                    <SPLIT distance="250" swimtime="00:04:18.79" />
                    <SPLIT distance="300" swimtime="00:05:14.40" />
                    <SPLIT distance="350" swimtime="00:05:56.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="336" swimtime="00:11:36.98" resultid="7770" heatid="10634" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                    <SPLIT distance="100" swimtime="00:01:18.75" />
                    <SPLIT distance="150" swimtime="00:02:02.53" />
                    <SPLIT distance="200" swimtime="00:02:47.02" />
                    <SPLIT distance="250" swimtime="00:03:31.22" />
                    <SPLIT distance="300" swimtime="00:04:15.44" />
                    <SPLIT distance="350" swimtime="00:04:59.29" />
                    <SPLIT distance="400" swimtime="00:05:43.90" />
                    <SPLIT distance="450" swimtime="00:06:27.91" />
                    <SPLIT distance="500" swimtime="00:07:13.14" />
                    <SPLIT distance="550" swimtime="00:07:57.63" />
                    <SPLIT distance="600" swimtime="00:08:42.00" />
                    <SPLIT distance="650" swimtime="00:09:26.38" />
                    <SPLIT distance="700" swimtime="00:10:10.61" />
                    <SPLIT distance="750" swimtime="00:10:54.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="381" swimtime="00:02:34.80" resultid="7771" heatid="10656" lane="6" entrytime="00:02:32.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                    <SPLIT distance="100" swimtime="00:01:15.42" />
                    <SPLIT distance="150" swimtime="00:01:56.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="359" swimtime="00:05:31.02" resultid="7772" heatid="10712" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                    <SPLIT distance="100" swimtime="00:01:16.07" />
                    <SPLIT distance="150" swimtime="00:01:58.49" />
                    <SPLIT distance="200" swimtime="00:02:40.87" />
                    <SPLIT distance="250" swimtime="00:03:24.18" />
                    <SPLIT distance="300" swimtime="00:04:07.32" />
                    <SPLIT distance="350" swimtime="00:04:50.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="309" swimtime="00:01:24.46" resultid="7773" heatid="10729" lane="2" entrytime="00:01:23.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Tolentino Smarczewski" birthdate="2008-09-01" gender="M" nation="BRA" license="378818" swrid="5596941" athleteid="7676" externalid="378818">
              <RESULTS>
                <RESULT eventid="1123" points="369" swimtime="00:10:30.26" resultid="7677" heatid="10514" lane="6" entrytime="00:09:41.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                    <SPLIT distance="100" swimtime="00:01:07.22" />
                    <SPLIT distance="150" swimtime="00:01:44.56" />
                    <SPLIT distance="200" swimtime="00:02:22.48" />
                    <SPLIT distance="250" swimtime="00:03:01.44" />
                    <SPLIT distance="300" swimtime="00:03:42.03" />
                    <SPLIT distance="350" swimtime="00:04:22.23" />
                    <SPLIT distance="400" swimtime="00:05:02.79" />
                    <SPLIT distance="450" swimtime="00:05:43.78" />
                    <SPLIT distance="500" swimtime="00:06:25.03" />
                    <SPLIT distance="550" swimtime="00:07:04.97" />
                    <SPLIT distance="600" swimtime="00:07:46.52" />
                    <SPLIT distance="650" swimtime="00:08:28.16" />
                    <SPLIT distance="700" swimtime="00:09:09.28" />
                    <SPLIT distance="750" swimtime="00:09:51.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="407" swimtime="00:02:49.19" resultid="7678" heatid="10491" lane="3" entrytime="00:02:46.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.57" />
                    <SPLIT distance="100" swimtime="00:01:19.95" />
                    <SPLIT distance="150" swimtime="00:02:03.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="373" swimtime="00:05:36.67" resultid="7679" heatid="10521" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.26" />
                    <SPLIT distance="100" swimtime="00:01:20.04" />
                    <SPLIT distance="150" swimtime="00:02:07.71" />
                    <SPLIT distance="200" swimtime="00:02:52.01" />
                    <SPLIT distance="250" swimtime="00:03:37.06" />
                    <SPLIT distance="300" swimtime="00:04:23.78" />
                    <SPLIT distance="350" swimtime="00:05:01.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="375" swimtime="00:01:18.83" resultid="7680" heatid="10597" lane="1" entrytime="00:01:17.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="442" swimtime="00:02:13.90" resultid="7681" heatid="10672" lane="6" entrytime="00:02:09.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                    <SPLIT distance="100" swimtime="00:01:03.90" />
                    <SPLIT distance="150" swimtime="00:01:39.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="382" swimtime="00:05:03.05" resultid="7682" heatid="10722" lane="7" entrytime="00:04:47.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                    <SPLIT distance="100" swimtime="00:01:10.14" />
                    <SPLIT distance="150" swimtime="00:01:48.44" />
                    <SPLIT distance="200" swimtime="00:02:27.77" />
                    <SPLIT distance="250" swimtime="00:03:08.04" />
                    <SPLIT distance="300" swimtime="00:03:48.19" />
                    <SPLIT distance="350" swimtime="00:04:25.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Do Prado Martins" birthdate="2008-10-17" gender="F" nation="BRA" license="369419" swrid="5596893" athleteid="7641" externalid="369419">
              <RESULTS>
                <RESULT eventid="1079" points="440" swimtime="00:03:00.80" resultid="7642" heatid="10486" lane="1" entrytime="00:02:54.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                    <SPLIT distance="100" swimtime="00:01:24.33" />
                    <SPLIT distance="150" swimtime="00:02:12.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="479" swimtime="00:00:37.26" resultid="7643" heatid="10565" lane="1" entrytime="00:00:36.69" entrycourse="LCM" />
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 16:56)" eventid="1131" status="DSQ" swimtime="00:05:40.21" resultid="7644" heatid="10520" lane="5" entrytime="00:05:35.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.03" />
                    <SPLIT distance="100" swimtime="00:01:12.69" />
                    <SPLIT distance="150" swimtime="00:01:57.32" />
                    <SPLIT distance="200" swimtime="00:02:41.52" />
                    <SPLIT distance="250" swimtime="00:03:29.64" />
                    <SPLIT distance="300" swimtime="00:04:19.17" />
                    <SPLIT distance="350" swimtime="00:05:00.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="457" swimtime="00:01:23.21" resultid="7645" heatid="10588" lane="5" entrytime="00:01:20.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="483" swimtime="00:02:40.72" resultid="7646" heatid="10644" lane="3" entrytime="00:02:35.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.22" />
                    <SPLIT distance="100" swimtime="00:01:17.13" />
                    <SPLIT distance="150" swimtime="00:02:04.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="456" swimtime="00:01:11.64" resultid="7647" heatid="10702" lane="6" entrytime="00:01:11.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hendrik" lastname="Alteiro Groenwold" birthdate="2011-03-23" gender="M" nation="BRA" license="365756" swrid="5588520" athleteid="7627" externalid="365756">
              <RESULTS>
                <RESULT eventid="1071" points="523" swimtime="00:02:18.84" resultid="7628" heatid="10480" lane="7" entrytime="00:02:19.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                    <SPLIT distance="100" swimtime="00:01:06.90" />
                    <SPLIT distance="150" swimtime="00:01:43.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="394" swimtime="00:02:30.42" resultid="7629" heatid="10558" lane="1" entrytime="00:02:23.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                    <SPLIT distance="100" swimtime="00:01:09.27" />
                    <SPLIT distance="150" swimtime="00:01:50.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="472" swimtime="00:18:38.18" resultid="7630" heatid="10638" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                    <SPLIT distance="100" swimtime="00:01:08.82" />
                    <SPLIT distance="150" swimtime="00:01:45.84" />
                    <SPLIT distance="200" swimtime="00:02:23.09" />
                    <SPLIT distance="250" swimtime="00:03:00.48" />
                    <SPLIT distance="300" swimtime="00:03:37.04" />
                    <SPLIT distance="350" swimtime="00:04:13.96" />
                    <SPLIT distance="400" swimtime="00:04:51.44" />
                    <SPLIT distance="450" swimtime="00:05:28.59" />
                    <SPLIT distance="500" swimtime="00:06:05.45" />
                    <SPLIT distance="550" swimtime="00:06:42.94" />
                    <SPLIT distance="600" swimtime="00:07:19.85" />
                    <SPLIT distance="650" swimtime="00:07:57.91" />
                    <SPLIT distance="700" swimtime="00:08:35.25" />
                    <SPLIT distance="750" swimtime="00:09:12.67" />
                    <SPLIT distance="800" swimtime="00:09:50.22" />
                    <SPLIT distance="850" swimtime="00:10:27.47" />
                    <SPLIT distance="900" swimtime="00:11:04.72" />
                    <SPLIT distance="950" swimtime="00:11:42.92" />
                    <SPLIT distance="1000" swimtime="00:12:20.33" />
                    <SPLIT distance="1050" swimtime="00:12:57.69" />
                    <SPLIT distance="1100" swimtime="00:13:35.91" />
                    <SPLIT distance="1150" swimtime="00:14:13.91" />
                    <SPLIT distance="1200" swimtime="00:14:52.35" />
                    <SPLIT distance="1250" swimtime="00:15:30.09" />
                    <SPLIT distance="1300" swimtime="00:16:07.83" />
                    <SPLIT distance="1350" swimtime="00:16:46.61" />
                    <SPLIT distance="1400" swimtime="00:17:24.34" />
                    <SPLIT distance="1450" swimtime="00:18:01.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="523" swimtime="00:02:06.52" resultid="7631" heatid="10672" lane="1" entrytime="00:02:09.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                    <SPLIT distance="100" swimtime="00:01:01.24" />
                    <SPLIT distance="150" swimtime="00:01:34.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="420" swimtime="00:01:05.98" resultid="7632" heatid="10710" lane="9" entrytime="00:01:04.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="499" swimtime="00:01:05.02" resultid="7633" heatid="10741" lane="6" entrytime="00:01:04.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Macedo Medeiros" birthdate="2012-05-12" gender="M" nation="BRA" license="392015" swrid="4697574" athleteid="7753" externalid="392015">
              <RESULTS>
                <RESULT eventid="1087" points="252" swimtime="00:03:18.61" resultid="7754" heatid="10487" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.99" />
                    <SPLIT distance="100" swimtime="00:01:35.44" />
                    <SPLIT distance="150" swimtime="00:02:28.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="218" swimtime="00:00:43.08" resultid="7755" heatid="10571" lane="0" entrytime="00:00:44.72" entrycourse="LCM" />
                <RESULT eventid="1219" points="236" swimtime="00:01:31.93" resultid="7756" heatid="10592" lane="7" entrytime="00:01:42.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="243" swimtime="00:03:02.46" resultid="7757" heatid="10646" lane="1" entrytime="00:03:21.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.36" />
                    <SPLIT distance="100" swimtime="00:01:32.13" />
                    <SPLIT distance="150" swimtime="00:02:22.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="151" swimtime="00:01:32.75" resultid="7758" heatid="10704" lane="4" entrytime="00:01:47.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="160" swimtime="00:01:34.97" resultid="7759" heatid="10734" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Breno" lastname="Zanella Janke" birthdate="2011-04-26" gender="M" nation="BRA" license="365697" swrid="5588970" athleteid="7648" externalid="365697">
              <RESULTS>
                <RESULT eventid="1123" points="447" swimtime="00:09:50.95" resultid="7649" heatid="10514" lane="7" entrytime="00:09:53.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                    <SPLIT distance="100" swimtime="00:01:06.92" />
                    <SPLIT distance="150" swimtime="00:01:44.07" />
                    <SPLIT distance="200" swimtime="00:02:20.14" />
                    <SPLIT distance="250" swimtime="00:02:56.49" />
                    <SPLIT distance="300" swimtime="00:03:33.57" />
                    <SPLIT distance="350" swimtime="00:04:10.90" />
                    <SPLIT distance="400" swimtime="00:04:47.93" />
                    <SPLIT distance="450" swimtime="00:05:25.89" />
                    <SPLIT distance="500" swimtime="00:06:04.54" />
                    <SPLIT distance="550" swimtime="00:06:43.19" />
                    <SPLIT distance="600" swimtime="00:07:22.19" />
                    <SPLIT distance="650" swimtime="00:07:59.87" />
                    <SPLIT distance="700" swimtime="00:08:38.62" />
                    <SPLIT distance="750" swimtime="00:09:14.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="357" swimtime="00:02:56.77" resultid="7650" heatid="10490" lane="3" entrytime="00:02:55.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.58" />
                    <SPLIT distance="100" swimtime="00:01:22.72" />
                    <SPLIT distance="150" swimtime="00:02:10.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="411" swimtime="00:05:26.11" resultid="7651" heatid="10522" lane="7" entrytime="00:05:21.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                    <SPLIT distance="100" swimtime="00:01:12.16" />
                    <SPLIT distance="150" swimtime="00:01:54.67" />
                    <SPLIT distance="200" swimtime="00:02:35.52" />
                    <SPLIT distance="250" swimtime="00:03:22.93" />
                    <SPLIT distance="300" swimtime="00:04:10.86" />
                    <SPLIT distance="350" swimtime="00:04:48.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="344" swimtime="00:01:21.11" resultid="7652" heatid="10595" lane="4" entrytime="00:01:20.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="427" swimtime="00:02:31.28" resultid="7653" heatid="10650" lane="4" entrytime="00:02:30.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                    <SPLIT distance="100" swimtime="00:01:09.66" />
                    <SPLIT distance="150" swimtime="00:01:57.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="450" swimtime="00:04:47.00" resultid="7654" heatid="10722" lane="8" entrytime="00:04:48.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                    <SPLIT distance="100" swimtime="00:01:07.09" />
                    <SPLIT distance="150" swimtime="00:01:44.59" />
                    <SPLIT distance="200" swimtime="00:02:21.32" />
                    <SPLIT distance="250" swimtime="00:02:59.98" />
                    <SPLIT distance="300" swimtime="00:03:38.88" />
                    <SPLIT distance="350" swimtime="00:04:13.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="Bortoli Da Silva" birthdate="2010-09-30" gender="M" nation="BRA" license="365500" swrid="4675666" athleteid="7774" externalid="365500">
              <RESULTS>
                <RESULT eventid="1103" points="367" swimtime="00:00:31.09" resultid="7775" heatid="10504" lane="3" entrytime="00:00:33.37" entrycourse="LCM" />
                <RESULT eventid="1171" points="352" swimtime="00:02:36.25" resultid="7776" heatid="10555" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                    <SPLIT distance="100" swimtime="00:01:13.29" />
                    <SPLIT distance="150" swimtime="00:01:55.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="400" swimtime="00:05:28.96" resultid="7777" heatid="10522" lane="9" entrytime="00:05:41.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                    <SPLIT distance="100" swimtime="00:01:11.14" />
                    <SPLIT distance="150" swimtime="00:01:56.04" />
                    <SPLIT distance="200" swimtime="00:02:40.81" />
                    <SPLIT distance="250" swimtime="00:03:27.74" />
                    <SPLIT distance="300" swimtime="00:04:16.93" />
                    <SPLIT distance="350" swimtime="00:04:54.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="397" swimtime="00:02:18.76" resultid="7778" heatid="10662" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                    <SPLIT distance="100" swimtime="00:01:06.72" />
                    <SPLIT distance="150" swimtime="00:01:42.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="352" swimtime="00:01:09.97" resultid="7779" heatid="10707" lane="2" entrytime="00:01:13.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="407" swimtime="00:04:56.82" resultid="7780" heatid="10718" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                    <SPLIT distance="100" swimtime="00:01:09.25" />
                    <SPLIT distance="150" swimtime="00:01:46.99" />
                    <SPLIT distance="200" swimtime="00:02:25.85" />
                    <SPLIT distance="250" swimtime="00:03:04.22" />
                    <SPLIT distance="300" swimtime="00:03:43.04" />
                    <SPLIT distance="350" swimtime="00:04:21.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Ramirez Vasconcelos" birthdate="2011-04-06" gender="M" nation="BRA" license="392013" swrid="4863662" athleteid="7746" externalid="392013">
              <RESULTS>
                <RESULT eventid="1087" points="452" swimtime="00:02:43.45" resultid="7747" heatid="10490" lane="5" entrytime="00:02:54.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="100" swimtime="00:01:17.07" />
                    <SPLIT distance="150" swimtime="00:02:00.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="362" swimtime="00:01:05.06" resultid="7748" heatid="10535" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="383" swimtime="00:05:33.80" resultid="7749" heatid="10521" lane="4" entrytime="00:05:52.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                    <SPLIT distance="100" swimtime="00:01:16.31" />
                    <SPLIT distance="150" swimtime="00:02:01.05" />
                    <SPLIT distance="200" swimtime="00:02:45.19" />
                    <SPLIT distance="250" swimtime="00:03:30.57" />
                    <SPLIT distance="300" swimtime="00:04:17.27" />
                    <SPLIT distance="350" swimtime="00:04:56.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="417" swimtime="00:01:16.11" resultid="7750" heatid="10595" lane="3" entrytime="00:01:21.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="413" swimtime="00:02:33.03" resultid="7751" heatid="10649" lane="8" entrytime="00:02:43.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                    <SPLIT distance="100" swimtime="00:01:14.19" />
                    <SPLIT distance="150" swimtime="00:01:56.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="329" swimtime="00:01:11.62" resultid="7752" heatid="10704" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Flavia" lastname="De Metz" birthdate="2011-01-07" gender="F" nation="BRA" license="390846" swrid="5596887" athleteid="7739" externalid="390846">
              <RESULTS>
                <RESULT eventid="1115" points="353" swimtime="00:21:42.42" resultid="7740" heatid="10512" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                    <SPLIT distance="100" swimtime="00:01:15.13" />
                    <SPLIT distance="150" swimtime="00:01:56.67" />
                    <SPLIT distance="200" swimtime="00:02:38.54" />
                    <SPLIT distance="250" swimtime="00:03:20.69" />
                    <SPLIT distance="300" swimtime="00:04:04.38" />
                    <SPLIT distance="350" swimtime="00:04:47.55" />
                    <SPLIT distance="400" swimtime="00:05:31.52" />
                    <SPLIT distance="450" swimtime="00:06:15.63" />
                    <SPLIT distance="500" swimtime="00:07:00.49" />
                    <SPLIT distance="550" swimtime="00:07:46.26" />
                    <SPLIT distance="600" swimtime="00:08:31.32" />
                    <SPLIT distance="650" swimtime="00:09:17.31" />
                    <SPLIT distance="700" swimtime="00:10:02.69" />
                    <SPLIT distance="750" swimtime="00:10:48.01" />
                    <SPLIT distance="800" swimtime="00:11:34.12" />
                    <SPLIT distance="850" swimtime="00:12:19.78" />
                    <SPLIT distance="900" swimtime="00:13:02.93" />
                    <SPLIT distance="950" swimtime="00:13:46.90" />
                    <SPLIT distance="1000" swimtime="00:14:31.11" />
                    <SPLIT distance="1050" swimtime="00:15:16.25" />
                    <SPLIT distance="1100" swimtime="00:16:00.63" />
                    <SPLIT distance="1150" swimtime="00:16:45.45" />
                    <SPLIT distance="1200" swimtime="00:17:28.91" />
                    <SPLIT distance="1250" swimtime="00:18:12.49" />
                    <SPLIT distance="1300" swimtime="00:18:55.13" />
                    <SPLIT distance="1350" swimtime="00:19:38.03" />
                    <SPLIT distance="1400" swimtime="00:20:20.16" />
                    <SPLIT distance="1450" swimtime="00:21:02.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="365" swimtime="00:02:52.30" resultid="7741" heatid="10471" lane="6" entrytime="00:02:52.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.76" />
                    <SPLIT distance="100" swimtime="00:01:23.46" />
                    <SPLIT distance="150" swimtime="00:02:09.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="474" swimtime="00:01:06.32" resultid="7742" heatid="10532" lane="0" entrytime="00:01:06.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="368" swimtime="00:11:16.29" resultid="7743" heatid="10632" lane="8" entrytime="00:10:45.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                    <SPLIT distance="100" swimtime="00:01:11.95" />
                    <SPLIT distance="150" swimtime="00:01:53.48" />
                    <SPLIT distance="200" swimtime="00:02:34.92" />
                    <SPLIT distance="250" swimtime="00:03:18.20" />
                    <SPLIT distance="300" swimtime="00:04:01.63" />
                    <SPLIT distance="350" swimtime="00:04:46.25" />
                    <SPLIT distance="400" swimtime="00:05:29.72" />
                    <SPLIT distance="450" swimtime="00:06:14.16" />
                    <SPLIT distance="500" swimtime="00:06:58.25" />
                    <SPLIT distance="550" swimtime="00:07:42.46" />
                    <SPLIT distance="600" swimtime="00:08:27.41" />
                    <SPLIT distance="650" swimtime="00:09:11.73" />
                    <SPLIT distance="700" swimtime="00:09:55.53" />
                    <SPLIT distance="750" swimtime="00:10:36.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="464" swimtime="00:02:24.87" resultid="7744" heatid="10658" lane="5" entrytime="00:02:24.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                    <SPLIT distance="100" swimtime="00:01:08.73" />
                    <SPLIT distance="150" swimtime="00:01:46.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="378" swimtime="00:05:25.36" resultid="7745" heatid="10715" lane="9" entrytime="00:05:11.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:13.35" />
                    <SPLIT distance="150" swimtime="00:01:55.59" />
                    <SPLIT distance="200" swimtime="00:02:37.00" />
                    <SPLIT distance="250" swimtime="00:03:20.43" />
                    <SPLIT distance="300" swimtime="00:04:03.67" />
                    <SPLIT distance="350" swimtime="00:04:46.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luann" lastname="Miguel Mazur" birthdate="2007-01-10" gender="M" nation="BRA" license="365682" swrid="5596915" athleteid="7620" externalid="365682">
              <RESULTS>
                <RESULT eventid="1087" points="385" swimtime="00:02:52.40" resultid="7621" heatid="10492" lane="9" entrytime="00:02:39.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.00" />
                    <SPLIT distance="100" swimtime="00:01:20.14" />
                    <SPLIT distance="150" swimtime="00:02:05.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="451" swimtime="00:00:33.83" resultid="7622" heatid="10574" lane="7" entrytime="00:00:34.21" entrycourse="LCM" />
                <RESULT comment="SW 6.4 - Não começou a executar a virada imediatamente após virar para a posição de peito.  (Horário: 17:17)" eventid="1139" status="DSQ" swimtime="00:05:37.72" resultid="7623" heatid="10523" lane="8" entrytime="00:05:07.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                    <SPLIT distance="100" swimtime="00:01:12.93" />
                    <SPLIT distance="150" swimtime="00:01:58.38" />
                    <SPLIT distance="200" swimtime="00:02:41.85" />
                    <SPLIT distance="250" swimtime="00:03:29.52" />
                    <SPLIT distance="300" swimtime="00:04:15.90" />
                    <SPLIT distance="350" swimtime="00:04:57.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="403" swimtime="00:01:16.95" resultid="7624" heatid="10597" lane="5" entrytime="00:01:14.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="365" swimtime="00:02:39.42" resultid="7625" heatid="10651" lane="7" entrytime="00:02:25.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                    <SPLIT distance="100" swimtime="00:01:16.15" />
                    <SPLIT distance="150" swimtime="00:02:02.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="336" swimtime="00:05:16.42" resultid="7626" heatid="10717" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                    <SPLIT distance="100" swimtime="00:01:13.87" />
                    <SPLIT distance="150" swimtime="00:01:54.05" />
                    <SPLIT distance="200" swimtime="00:02:35.28" />
                    <SPLIT distance="250" swimtime="00:03:16.92" />
                    <SPLIT distance="300" swimtime="00:03:58.95" />
                    <SPLIT distance="350" swimtime="00:04:37.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Claudio" lastname="Rohnelt" birthdate="2010-03-08" gender="M" nation="BRA" license="357954" swrid="5596935" athleteid="7613" externalid="357954">
              <RESULTS>
                <RESULT eventid="1123" points="344" swimtime="00:10:45.19" resultid="7614" heatid="10515" lane="1" entrytime="00:10:22.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                    <SPLIT distance="100" swimtime="00:01:11.79" />
                    <SPLIT distance="150" swimtime="00:01:51.11" />
                    <SPLIT distance="200" swimtime="00:02:31.53" />
                    <SPLIT distance="250" swimtime="00:03:11.53" />
                    <SPLIT distance="300" swimtime="00:03:52.16" />
                    <SPLIT distance="350" swimtime="00:04:32.91" />
                    <SPLIT distance="400" swimtime="00:05:13.82" />
                    <SPLIT distance="450" swimtime="00:05:55.06" />
                    <SPLIT distance="500" swimtime="00:06:36.11" />
                    <SPLIT distance="550" swimtime="00:07:17.81" />
                    <SPLIT distance="600" swimtime="00:07:59.24" />
                    <SPLIT distance="650" swimtime="00:08:40.49" />
                    <SPLIT distance="700" swimtime="00:09:21.68" />
                    <SPLIT distance="750" swimtime="00:10:03.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="298" swimtime="00:02:45.02" resultid="7615" heatid="10556" lane="5" entrytime="00:02:41.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="100" swimtime="00:01:14.56" />
                    <SPLIT distance="150" swimtime="00:01:58.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="346" swimtime="00:20:39.69" resultid="7616" heatid="10637" lane="1" entrytime="00:20:46.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                    <SPLIT distance="100" swimtime="00:01:13.89" />
                    <SPLIT distance="150" swimtime="00:01:53.73" />
                    <SPLIT distance="200" swimtime="00:02:33.92" />
                    <SPLIT distance="250" swimtime="00:03:14.14" />
                    <SPLIT distance="300" swimtime="00:03:54.53" />
                    <SPLIT distance="350" swimtime="00:04:34.71" />
                    <SPLIT distance="400" swimtime="00:05:15.43" />
                    <SPLIT distance="450" swimtime="00:05:56.34" />
                    <SPLIT distance="500" swimtime="00:06:37.45" />
                    <SPLIT distance="550" swimtime="00:07:18.73" />
                    <SPLIT distance="600" swimtime="00:08:00.48" />
                    <SPLIT distance="650" swimtime="00:08:41.80" />
                    <SPLIT distance="700" swimtime="00:09:23.14" />
                    <SPLIT distance="750" swimtime="00:10:04.88" />
                    <SPLIT distance="800" swimtime="00:10:46.88" />
                    <SPLIT distance="850" swimtime="00:11:29.03" />
                    <SPLIT distance="900" swimtime="00:12:11.00" />
                    <SPLIT distance="950" swimtime="00:12:53.11" />
                    <SPLIT distance="1000" swimtime="00:13:36.17" />
                    <SPLIT distance="1050" swimtime="00:14:18.19" />
                    <SPLIT distance="1100" swimtime="00:15:01.02" />
                    <SPLIT distance="1150" swimtime="00:15:43.40" />
                    <SPLIT distance="1200" swimtime="00:16:26.05" />
                    <SPLIT distance="1250" swimtime="00:17:08.94" />
                    <SPLIT distance="1300" swimtime="00:17:51.41" />
                    <SPLIT distance="1350" swimtime="00:18:33.77" />
                    <SPLIT distance="1400" swimtime="00:19:16.14" />
                    <SPLIT distance="1450" swimtime="00:19:58.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="363" swimtime="00:02:39.73" resultid="7617" heatid="10645" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                    <SPLIT distance="100" swimtime="00:01:14.07" />
                    <SPLIT distance="150" swimtime="00:02:02.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="269" swimtime="00:01:16.54" resultid="7618" heatid="10707" lane="5" entrytime="00:01:12.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="369" swimtime="00:05:06.65" resultid="7619" heatid="10720" lane="2" entrytime="00:05:10.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                    <SPLIT distance="100" swimtime="00:01:10.95" />
                    <SPLIT distance="150" swimtime="00:01:50.05" />
                    <SPLIT distance="200" swimtime="00:02:29.22" />
                    <SPLIT distance="250" swimtime="00:03:08.51" />
                    <SPLIT distance="300" swimtime="00:03:47.72" />
                    <SPLIT distance="350" swimtime="00:04:27.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="16" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1205" points="538" swimtime="00:08:34.60" resultid="7807" heatid="10580" lane="3" entrytime="00:08:27.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.50" />
                    <SPLIT distance="100" swimtime="00:01:02.58" />
                    <SPLIT distance="150" swimtime="00:01:36.95" />
                    <SPLIT distance="200" swimtime="00:02:11.11" />
                    <SPLIT distance="250" swimtime="00:02:40.90" />
                    <SPLIT distance="300" swimtime="00:03:13.77" />
                    <SPLIT distance="350" swimtime="00:03:47.83" />
                    <SPLIT distance="400" swimtime="00:04:20.80" />
                    <SPLIT distance="450" swimtime="00:04:50.03" />
                    <SPLIT distance="500" swimtime="00:05:21.97" />
                    <SPLIT distance="550" swimtime="00:05:55.09" />
                    <SPLIT distance="600" swimtime="00:06:28.05" />
                    <SPLIT distance="650" swimtime="00:06:56.18" />
                    <SPLIT distance="700" swimtime="00:07:27.89" />
                    <SPLIT distance="750" swimtime="00:08:01.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7704" number="1" />
                    <RELAYPOSITION athleteid="7669" number="2" />
                    <RELAYPOSITION athleteid="7585" number="3" />
                    <RELAYPOSITION athleteid="7606" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="19" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1207" points="521" swimtime="00:08:39.96" resultid="7808" heatid="10581" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.05" />
                    <SPLIT distance="100" swimtime="00:00:59.79" />
                    <SPLIT distance="150" swimtime="00:01:33.94" />
                    <SPLIT distance="200" swimtime="00:02:08.37" />
                    <SPLIT distance="250" swimtime="00:02:37.49" />
                    <SPLIT distance="300" swimtime="00:03:10.43" />
                    <SPLIT distance="350" swimtime="00:03:45.30" />
                    <SPLIT distance="400" swimtime="00:04:20.07" />
                    <SPLIT distance="450" swimtime="00:04:49.90" />
                    <SPLIT distance="500" swimtime="00:05:23.26" />
                    <SPLIT distance="550" swimtime="00:05:59.12" />
                    <SPLIT distance="600" swimtime="00:06:37.14" />
                    <SPLIT distance="650" swimtime="00:07:04.66" />
                    <SPLIT distance="700" swimtime="00:07:35.75" />
                    <SPLIT distance="750" swimtime="00:08:07.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7711" number="1" />
                    <RELAYPOSITION athleteid="7676" number="2" />
                    <RELAYPOSITION athleteid="7620" number="3" />
                    <RELAYPOSITION athleteid="7571" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1203" points="450" swimtime="00:09:06.18" resultid="7809" heatid="10579" lane="5" entrytime="00:09:19.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.08" />
                    <SPLIT distance="100" swimtime="00:01:03.52" />
                    <SPLIT distance="150" swimtime="00:01:38.50" />
                    <SPLIT distance="200" swimtime="00:02:13.86" />
                    <SPLIT distance="250" swimtime="00:02:44.87" />
                    <SPLIT distance="300" swimtime="00:03:20.47" />
                    <SPLIT distance="350" swimtime="00:03:57.28" />
                    <SPLIT distance="400" swimtime="00:04:33.05" />
                    <SPLIT distance="450" swimtime="00:05:04.81" />
                    <SPLIT distance="500" swimtime="00:05:41.43" />
                    <SPLIT distance="550" swimtime="00:06:19.40" />
                    <SPLIT distance="600" swimtime="00:06:56.01" />
                    <SPLIT distance="650" swimtime="00:07:23.90" />
                    <SPLIT distance="700" swimtime="00:07:56.42" />
                    <SPLIT distance="750" swimtime="00:08:31.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7648" number="1" />
                    <RELAYPOSITION athleteid="7746" number="2" />
                    <RELAYPOSITION athleteid="7662" number="3" />
                    <RELAYPOSITION athleteid="7627" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1331" points="496" swimtime="00:04:21.06" resultid="7810" heatid="10698" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                    <SPLIT distance="100" swimtime="00:01:07.20" />
                    <SPLIT distance="150" swimtime="00:01:42.44" />
                    <SPLIT distance="200" swimtime="00:02:23.81" />
                    <SPLIT distance="250" swimtime="00:02:53.59" />
                    <SPLIT distance="300" swimtime="00:03:26.41" />
                    <SPLIT distance="350" swimtime="00:03:52.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7795" number="1" />
                    <RELAYPOSITION athleteid="7676" number="2" />
                    <RELAYPOSITION athleteid="7711" number="3" />
                    <RELAYPOSITION athleteid="7571" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1399" points="510" swimtime="00:03:55.52" resultid="7813" heatid="10753" lane="1" entrytime="00:04:06.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.09" />
                    <SPLIT distance="100" swimtime="00:00:55.76" />
                    <SPLIT distance="150" swimtime="00:01:23.89" />
                    <SPLIT distance="200" swimtime="00:01:55.59" />
                    <SPLIT distance="250" swimtime="00:02:23.63" />
                    <SPLIT distance="300" swimtime="00:02:56.50" />
                    <SPLIT distance="350" swimtime="00:03:24.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7571" number="1" />
                    <RELAYPOSITION athleteid="7711" number="2" />
                    <RELAYPOSITION athleteid="7795" number="3" />
                    <RELAYPOSITION athleteid="7676" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1327" points="421" swimtime="00:04:35.83" resultid="7811" heatid="10696" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                    <SPLIT distance="100" swimtime="00:01:07.39" />
                    <SPLIT distance="150" swimtime="00:01:44.90" />
                    <SPLIT distance="200" swimtime="00:02:25.83" />
                    <SPLIT distance="250" swimtime="00:02:58.07" />
                    <SPLIT distance="300" swimtime="00:03:34.55" />
                    <SPLIT distance="350" swimtime="00:04:03.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7704" number="1" />
                    <RELAYPOSITION athleteid="7606" number="2" />
                    <RELAYPOSITION athleteid="7774" number="3" />
                    <RELAYPOSITION athleteid="7613" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1395" points="459" swimtime="00:04:03.99" resultid="7814" heatid="10751" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.20" />
                    <SPLIT distance="100" swimtime="00:01:00.42" />
                    <SPLIT distance="150" swimtime="00:01:29.84" />
                    <SPLIT distance="200" swimtime="00:02:02.81" />
                    <SPLIT distance="250" swimtime="00:02:33.37" />
                    <SPLIT distance="300" swimtime="00:03:06.71" />
                    <SPLIT distance="350" swimtime="00:03:34.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7704" number="1" />
                    <RELAYPOSITION athleteid="7613" number="2" />
                    <RELAYPOSITION athleteid="7774" number="3" />
                    <RELAYPOSITION athleteid="7606" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1325" points="459" swimtime="00:04:28.06" resultid="7812" heatid="10695" lane="6" entrytime="00:04:56.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                    <SPLIT distance="100" swimtime="00:01:04.79" />
                    <SPLIT distance="150" swimtime="00:01:40.13" />
                    <SPLIT distance="200" swimtime="00:02:21.02" />
                    <SPLIT distance="250" swimtime="00:02:52.13" />
                    <SPLIT distance="300" swimtime="00:03:26.64" />
                    <SPLIT distance="350" swimtime="00:03:55.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7627" number="1" />
                    <RELAYPOSITION athleteid="7746" number="2" />
                    <RELAYPOSITION athleteid="7648" number="3" />
                    <RELAYPOSITION athleteid="7725" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1393" points="455" swimtime="00:04:04.72" resultid="7815" heatid="10750" lane="3" entrytime="00:04:12.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                    <SPLIT distance="100" swimtime="00:00:59.90" />
                    <SPLIT distance="150" swimtime="00:01:29.66" />
                    <SPLIT distance="200" swimtime="00:02:02.08" />
                    <SPLIT distance="250" swimtime="00:02:32.16" />
                    <SPLIT distance="300" swimtime="00:03:05.28" />
                    <SPLIT distance="350" swimtime="00:03:33.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7648" number="1" />
                    <RELAYPOSITION athleteid="7725" number="2" />
                    <RELAYPOSITION athleteid="7746" number="3" />
                    <RELAYPOSITION athleteid="7627" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="COMERCIAL CASCAVEL &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1325" points="303" swimtime="00:05:07.53" resultid="7798" heatid="10695" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.94" />
                    <SPLIT distance="100" swimtime="00:01:24.89" />
                    <SPLIT distance="150" swimtime="00:02:03.27" />
                    <SPLIT distance="200" swimtime="00:02:47.74" />
                    <SPLIT distance="250" swimtime="00:03:20.50" />
                    <SPLIT distance="300" swimtime="00:03:59.05" />
                    <SPLIT distance="350" swimtime="00:04:31.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7634" number="1" />
                    <RELAYPOSITION athleteid="7683" number="2" />
                    <RELAYPOSITION athleteid="7662" number="3" />
                    <RELAYPOSITION athleteid="7781" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1393" points="318" swimtime="00:04:35.77" resultid="7799" heatid="10749" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.13" />
                    <SPLIT distance="100" swimtime="00:01:05.46" />
                    <SPLIT distance="150" swimtime="00:01:38.54" />
                    <SPLIT distance="200" swimtime="00:02:14.92" />
                    <SPLIT distance="250" swimtime="00:02:49.14" />
                    <SPLIT distance="300" swimtime="00:03:26.80" />
                    <SPLIT distance="350" swimtime="00:03:59.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7662" number="1" />
                    <RELAYPOSITION athleteid="7718" number="2" />
                    <RELAYPOSITION athleteid="7683" number="3" />
                    <RELAYPOSITION athleteid="7781" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="F" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1197" points="437" swimtime="00:10:02.69" resultid="7801" heatid="10577" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                    <SPLIT distance="100" swimtime="00:01:13.66" />
                    <SPLIT distance="150" swimtime="00:01:53.51" />
                    <SPLIT distance="200" swimtime="00:02:30.97" />
                    <SPLIT distance="250" swimtime="00:03:02.61" />
                    <SPLIT distance="300" swimtime="00:03:38.03" />
                    <SPLIT distance="350" swimtime="00:04:15.95" />
                    <SPLIT distance="400" swimtime="00:04:53.62" />
                    <SPLIT distance="450" swimtime="00:05:27.72" />
                    <SPLIT distance="500" swimtime="00:06:08.61" />
                    <SPLIT distance="550" swimtime="00:06:49.57" />
                    <SPLIT distance="600" swimtime="00:07:30.09" />
                    <SPLIT distance="650" swimtime="00:08:06.06" />
                    <SPLIT distance="750" swimtime="00:09:24.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7767" number="1" />
                    <RELAYPOSITION athleteid="7697" number="2" />
                    <RELAYPOSITION athleteid="7592" number="3" />
                    <RELAYPOSITION athleteid="7599" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1195" points="384" swimtime="00:10:29.08" resultid="7802" heatid="10576" lane="3" entrytime="00:09:58.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                    <SPLIT distance="100" swimtime="00:01:11.42" />
                    <SPLIT distance="150" swimtime="00:01:50.69" />
                    <SPLIT distance="200" swimtime="00:02:29.82" />
                    <SPLIT distance="250" swimtime="00:03:07.27" />
                    <SPLIT distance="300" swimtime="00:03:50.76" />
                    <SPLIT distance="350" swimtime="00:04:35.88" />
                    <SPLIT distance="500" swimtime="00:06:38.83" />
                    <SPLIT distance="550" swimtime="00:07:20.70" />
                    <SPLIT distance="650" swimtime="00:08:33.74" />
                    <SPLIT distance="700" swimtime="00:09:10.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7739" number="1" />
                    <RELAYPOSITION athleteid="7760" number="2" />
                    <RELAYPOSITION athleteid="7690" number="3" />
                    <RELAYPOSITION athleteid="7655" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1315" points="347" swimtime="00:05:26.54" resultid="7803" heatid="10689" lane="7" entrytime="00:05:03.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.37" />
                    <SPLIT distance="100" swimtime="00:01:22.17" />
                    <SPLIT distance="150" swimtime="00:02:03.90" />
                    <SPLIT distance="200" swimtime="00:02:50.82" />
                    <SPLIT distance="250" swimtime="00:03:30.07" />
                    <SPLIT distance="300" swimtime="00:04:17.78" />
                    <SPLIT distance="350" swimtime="00:04:50.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7739" number="1" />
                    <RELAYPOSITION athleteid="7690" number="2" />
                    <RELAYPOSITION athleteid="7760" number="3" />
                    <RELAYPOSITION athleteid="7655" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1383" points="371" swimtime="00:04:49.37" resultid="7806" heatid="10744" lane="5" entrytime="00:04:30.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.26" />
                    <SPLIT distance="100" swimtime="00:01:06.54" />
                    <SPLIT distance="150" swimtime="00:01:43.29" />
                    <SPLIT distance="200" swimtime="00:02:23.44" />
                    <SPLIT distance="250" swimtime="00:02:59.44" />
                    <SPLIT distance="300" swimtime="00:03:39.31" />
                    <SPLIT distance="350" swimtime="00:04:12.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7739" number="1" />
                    <RELAYPOSITION athleteid="7690" number="2" />
                    <RELAYPOSITION athleteid="7760" number="3" />
                    <RELAYPOSITION athleteid="7655" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="F" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1319" points="422" swimtime="00:05:06.09" resultid="7804" heatid="10691" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                    <SPLIT distance="100" swimtime="00:01:15.44" />
                    <SPLIT distance="150" swimtime="00:01:53.02" />
                    <SPLIT distance="200" swimtime="00:02:36.74" />
                    <SPLIT distance="250" swimtime="00:03:13.64" />
                    <SPLIT distance="300" swimtime="00:03:57.56" />
                    <SPLIT distance="350" swimtime="00:04:30.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7592" number="1" />
                    <RELAYPOSITION athleteid="7697" number="2" />
                    <RELAYPOSITION athleteid="7599" number="3" />
                    <RELAYPOSITION athleteid="7767" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1387" points="431" swimtime="00:04:35.23" resultid="7805" heatid="10746" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                    <SPLIT distance="100" swimtime="00:01:08.92" />
                    <SPLIT distance="150" swimtime="00:01:40.95" />
                    <SPLIT distance="200" swimtime="00:02:15.40" />
                    <SPLIT distance="250" swimtime="00:02:48.92" />
                    <SPLIT distance="300" swimtime="00:03:27.62" />
                    <SPLIT distance="350" swimtime="00:04:00.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7599" number="1" />
                    <RELAYPOSITION athleteid="7697" number="2" />
                    <RELAYPOSITION athleteid="7592" number="3" />
                    <RELAYPOSITION athleteid="7767" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1113" points="424" swimtime="00:04:49.36" resultid="7816" heatid="10510" lane="5" entrytime="00:04:51.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="100" swimtime="00:01:06.04" />
                    <SPLIT distance="150" swimtime="00:01:47.84" />
                    <SPLIT distance="200" swimtime="00:02:35.04" />
                    <SPLIT distance="250" swimtime="00:03:07.11" />
                    <SPLIT distance="300" swimtime="00:03:43.37" />
                    <SPLIT distance="350" swimtime="00:04:15.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7627" number="1" />
                    <RELAYPOSITION athleteid="7690" number="2" />
                    <RELAYPOSITION athleteid="7648" number="3" />
                    <RELAYPOSITION athleteid="7739" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="X" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1247" points="483" swimtime="00:04:36.94" resultid="7817" heatid="10631" lane="6" entrytime="00:04:45.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.08" />
                    <SPLIT distance="100" swimtime="00:01:03.91" />
                    <SPLIT distance="150" swimtime="00:01:42.98" />
                    <SPLIT distance="200" swimtime="00:02:27.47" />
                    <SPLIT distance="250" swimtime="00:02:57.00" />
                    <SPLIT distance="300" swimtime="00:03:28.95" />
                    <SPLIT distance="350" swimtime="00:04:01.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7571" number="1" />
                    <RELAYPOSITION athleteid="7641" number="2" />
                    <RELAYPOSITION athleteid="7711" number="3" />
                    <RELAYPOSITION athleteid="7564" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="X" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1243" points="459" swimtime="00:04:41.68" resultid="7818" heatid="10629" lane="2" entrytime="00:04:46.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="100" swimtime="00:01:14.67" />
                    <SPLIT distance="150" swimtime="00:01:53.88" />
                    <SPLIT distance="200" swimtime="00:02:37.21" />
                    <SPLIT distance="250" swimtime="00:03:09.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7592" number="1" />
                    <RELAYPOSITION athleteid="7697" number="2" />
                    <RELAYPOSITION athleteid="7704" number="3" />
                    <RELAYPOSITION athleteid="7606" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="X" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1245" points="458" swimtime="00:04:41.87" resultid="7819" heatid="10630" lane="3" entrytime="00:04:32.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                    <SPLIT distance="100" swimtime="00:01:16.01" />
                    <SPLIT distance="150" swimtime="00:01:51.40" />
                    <SPLIT distance="200" swimtime="00:02:32.48" />
                    <SPLIT distance="300" swimtime="00:03:33.44" />
                    <SPLIT distance="350" swimtime="00:04:05.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7599" number="1" />
                    <RELAYPOSITION athleteid="7585" number="2" />
                    <RELAYPOSITION athleteid="7669" number="3" />
                    <RELAYPOSITION athleteid="7767" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="COMERCIAL CASCAVEL &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1113" points="373" swimtime="00:05:01.83" resultid="7800" heatid="10510" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.76" />
                    <SPLIT distance="150" swimtime="00:01:59.82" />
                    <SPLIT distance="200" swimtime="00:02:41.61" />
                    <SPLIT distance="250" swimtime="00:03:14.62" />
                    <SPLIT distance="300" swimtime="00:03:52.61" />
                    <SPLIT distance="350" swimtime="00:04:25.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7760" number="1" />
                    <RELAYPOSITION athleteid="7746" number="2" />
                    <RELAYPOSITION athleteid="7662" number="3" />
                    <RELAYPOSITION athleteid="7655" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="19584" nation="BRA" region="SC" clubid="7260" name="Clube De Caca E Tiro Vasconcelos Drumond" shortname="Atiradores Natação">
          <ATHLETES>
            <ATHLETE firstname="Vinicius" lastname="Decker Ferrari" birthdate="2008-11-21" gender="M" nation="BRA" license="382021" swrid="5736534" athleteid="7267" externalid="382021">
              <RESULTS>
                <RESULT eventid="1155" points="529" status="EXH" swimtime="00:00:57.36" resultid="7268" heatid="10550" lane="6" entrytime="00:00:56.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="536" status="EXH" swimtime="00:00:25.74" resultid="7269" heatid="10626" lane="4" entrytime="00:00:25.54" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Ogata" birthdate="2010-01-06" gender="M" nation="BRA" license="388204" swrid="5634741" athleteid="7274" externalid="388204">
              <RESULTS>
                <RESULT eventid="1155" points="507" status="EXH" swimtime="00:00:58.18" resultid="7275" heatid="10547" lane="7" entrytime="00:01:01.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="451" status="EXH" swimtime="00:00:27.26" resultid="7276" heatid="10622" lane="9" entrytime="00:00:28.33" entrycourse="LCM" />
                <RESULT eventid="1273" points="429" status="EXH" swimtime="00:02:31.13" resultid="7277" heatid="10651" lane="8" entrytime="00:02:28.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                    <SPLIT distance="100" swimtime="00:01:11.95" />
                    <SPLIT distance="150" swimtime="00:01:56.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="528" status="EXH" swimtime="00:04:32.15" resultid="7278" heatid="10721" lane="1" entrytime="00:04:58.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                    <SPLIT distance="100" swimtime="00:01:04.34" />
                    <SPLIT distance="150" swimtime="00:01:39.04" />
                    <SPLIT distance="200" swimtime="00:02:13.85" />
                    <SPLIT distance="250" swimtime="00:02:48.67" />
                    <SPLIT distance="300" swimtime="00:03:23.71" />
                    <SPLIT distance="350" swimtime="00:03:58.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="José" lastname="Henrique Vargas Neto" birthdate="2007-06-29" gender="M" nation="BRA" license="353642" swrid="5736535" athleteid="7261" externalid="353642">
              <RESULTS>
                <RESULT eventid="1071" points="317" status="EXH" swimtime="00:02:43.98" resultid="7262" heatid="10477" lane="4" entrytime="00:02:36.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                    <SPLIT distance="100" swimtime="00:01:16.75" />
                    <SPLIT distance="150" swimtime="00:02:00.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="402" status="EXH" swimtime="00:01:02.86" resultid="7263" heatid="10548" lane="8" entrytime="00:01:00.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="408" status="EXH" swimtime="00:00:28.19" resultid="7264" heatid="10624" lane="1" entrytime="00:00:27.34" entrycourse="LCM" />
                <RESULT eventid="1305" points="447" status="EXH" swimtime="00:00:30.80" resultid="7265" heatid="10687" lane="1" entrytime="00:00:30.19" entrycourse="LCM" />
                <RESULT eventid="1373" points="401" status="EXH" swimtime="00:01:09.92" resultid="7266" heatid="10740" lane="0" entrytime="00:01:09.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Augusto" lastname="Mutz" birthdate="2009-04-23" gender="M" nation="BRA" license="382022" swrid="5634733" athleteid="7270" externalid="382022">
              <RESULTS>
                <RESULT eventid="1123" points="501" status="EXH" swimtime="00:09:28.92" resultid="7271" heatid="10514" lane="3" entrytime="00:09:38.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.53" />
                    <SPLIT distance="100" swimtime="00:01:05.58" />
                    <SPLIT distance="150" swimtime="00:01:40.58" />
                    <SPLIT distance="200" swimtime="00:02:15.91" />
                    <SPLIT distance="250" swimtime="00:02:51.61" />
                    <SPLIT distance="300" swimtime="00:03:27.30" />
                    <SPLIT distance="350" swimtime="00:04:03.47" />
                    <SPLIT distance="400" swimtime="00:04:39.38" />
                    <SPLIT distance="450" swimtime="00:05:15.38" />
                    <SPLIT distance="500" swimtime="00:05:51.52" />
                    <SPLIT distance="550" swimtime="00:06:27.93" />
                    <SPLIT distance="600" swimtime="00:07:04.18" />
                    <SPLIT distance="650" swimtime="00:07:40.89" />
                    <SPLIT distance="700" swimtime="00:08:17.18" />
                    <SPLIT distance="750" swimtime="00:08:53.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="512" status="EXH" swimtime="00:18:07.94" resultid="7272" heatid="10635" lane="8" entrytime="00:18:05.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                    <SPLIT distance="100" swimtime="00:01:07.38" />
                    <SPLIT distance="150" swimtime="00:01:43.40" />
                    <SPLIT distance="200" swimtime="00:02:19.46" />
                    <SPLIT distance="250" swimtime="00:02:55.72" />
                    <SPLIT distance="300" swimtime="00:03:32.25" />
                    <SPLIT distance="350" swimtime="00:04:09.03" />
                    <SPLIT distance="400" swimtime="00:04:45.55" />
                    <SPLIT distance="450" swimtime="00:05:21.49" />
                    <SPLIT distance="500" swimtime="00:05:58.09" />
                    <SPLIT distance="550" swimtime="00:06:34.67" />
                    <SPLIT distance="600" swimtime="00:07:11.05" />
                    <SPLIT distance="650" swimtime="00:07:47.67" />
                    <SPLIT distance="700" swimtime="00:08:24.11" />
                    <SPLIT distance="750" swimtime="00:09:00.20" />
                    <SPLIT distance="800" swimtime="00:09:36.83" />
                    <SPLIT distance="850" swimtime="00:10:13.48" />
                    <SPLIT distance="900" swimtime="00:10:50.11" />
                    <SPLIT distance="950" swimtime="00:11:26.96" />
                    <SPLIT distance="1000" swimtime="00:12:03.78" />
                    <SPLIT distance="1050" swimtime="00:12:40.53" />
                    <SPLIT distance="1100" swimtime="00:13:17.37" />
                    <SPLIT distance="1150" swimtime="00:13:54.00" />
                    <SPLIT distance="1200" swimtime="00:14:30.72" />
                    <SPLIT distance="1250" swimtime="00:15:07.42" />
                    <SPLIT distance="1300" swimtime="00:15:44.32" />
                    <SPLIT distance="1350" swimtime="00:16:21.47" />
                    <SPLIT distance="1400" swimtime="00:16:58.10" />
                    <SPLIT distance="1450" swimtime="00:17:33.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="505" status="EXH" swimtime="00:04:36.32" resultid="7273" heatid="10723" lane="2" entrytime="00:04:35.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.89" />
                    <SPLIT distance="100" swimtime="00:01:04.61" />
                    <SPLIT distance="150" swimtime="00:01:39.47" />
                    <SPLIT distance="200" swimtime="00:02:15.04" />
                    <SPLIT distance="250" swimtime="00:02:51.13" />
                    <SPLIT distance="300" swimtime="00:03:26.83" />
                    <SPLIT distance="350" swimtime="00:04:02.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="12782" nation="BRA" region="PR" clubid="8455" swrid="93773" name="Clube Duque De Caxias" shortname="Duque De Caxias">
          <ATHLETES>
            <ATHLETE firstname="Arthur" lastname="Gioia Brito" birthdate="2011-11-05" gender="M" nation="BRA" license="421525" swrid="5810757" athleteid="8499" externalid="421525">
              <RESULTS>
                <RESULT eventid="1087" points="261" swimtime="00:03:16.21" resultid="8500" heatid="10487" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.73" />
                    <SPLIT distance="100" swimtime="00:01:31.75" />
                    <SPLIT distance="150" swimtime="00:02:25.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="330" swimtime="00:00:37.52" resultid="8501" heatid="10568" lane="7" />
                <RESULT eventid="1235" points="323" swimtime="00:00:30.47" resultid="8502" heatid="10619" lane="1" entrytime="00:00:29.91" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ian" lastname="Berger" birthdate="2011-07-27" gender="M" nation="BRA" license="387966" swrid="5652879" athleteid="8469" externalid="387966">
              <RESULTS>
                <RESULT eventid="1103" points="293" swimtime="00:00:33.50" resultid="8470" heatid="10500" lane="6" />
                <RESULT eventid="1155" points="376" swimtime="00:01:04.24" resultid="8471" heatid="10545" lane="6" entrytime="00:01:04.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="366" swimtime="00:00:29.21" resultid="8472" heatid="10619" lane="3" entrytime="00:00:29.82" entrycourse="LCM" />
                <RESULT eventid="1357" points="360" swimtime="00:05:09.09" resultid="8473" heatid="10718" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                    <SPLIT distance="100" swimtime="00:01:10.97" />
                    <SPLIT distance="150" swimtime="00:01:49.73" />
                    <SPLIT distance="200" swimtime="00:02:29.21" />
                    <SPLIT distance="250" swimtime="00:03:08.83" />
                    <SPLIT distance="300" swimtime="00:03:49.10" />
                    <SPLIT distance="350" swimtime="00:04:29.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Flavia Braz" birthdate="2004-10-25" gender="F" nation="BRA" license="280573" swrid="5622281" athleteid="8456" externalid="280573">
              <RESULTS>
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="8457" heatid="10485" lane="7" entrytime="00:02:58.65" entrycourse="LCM" />
                <RESULT eventid="1179" points="546" swimtime="00:00:35.66" resultid="8458" heatid="10565" lane="6" entrytime="00:00:35.80" entrycourse="LCM" />
                <RESULT eventid="1211" points="493" swimtime="00:01:21.16" resultid="8459" heatid="10589" lane="3" entrytime="00:01:18.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="478" swimtime="00:02:23.50" resultid="8460" heatid="10653" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                    <SPLIT distance="100" swimtime="00:01:09.63" />
                    <SPLIT distance="150" swimtime="00:01:46.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" status="DNS" swimtime="00:00:00.00" resultid="8461" heatid="10699" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Kovalhuk Lima" birthdate="2009-03-16" gender="M" nation="BRA" license="417452" swrid="5762082" athleteid="8490" externalid="417452">
              <RESULTS>
                <RESULT eventid="1103" status="DNS" swimtime="00:00:00.00" resultid="8491" heatid="10501" lane="6" />
                <RESULT eventid="1155" points="369" swimtime="00:01:04.68" resultid="8492" heatid="10544" lane="4" entrytime="00:01:05.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="381" swimtime="00:00:28.84" resultid="8493" heatid="10610" lane="6" />
                <RESULT eventid="1305" points="299" swimtime="00:00:35.19" resultid="8494" heatid="10683" lane="9" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Vitor Girelli" birthdate="2009-08-01" gender="M" nation="BRA" license="387965" swrid="5622312" athleteid="8462" externalid="387965">
              <RESULTS>
                <RESULT eventid="1071" points="412" swimtime="00:02:30.40" resultid="8463" heatid="10474" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.71" />
                    <SPLIT distance="100" swimtime="00:01:11.96" />
                    <SPLIT distance="150" swimtime="00:01:51.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="317" swimtime="00:00:38.05" resultid="8464" heatid="10569" lane="6" />
                <RESULT eventid="1155" points="445" swimtime="00:01:00.77" resultid="8465" heatid="10547" lane="3" entrytime="00:01:01.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="401" swimtime="00:00:28.35" resultid="8466" heatid="10622" lane="2" entrytime="00:00:28.03" entrycourse="LCM" />
                <RESULT eventid="1305" points="384" swimtime="00:00:32.39" resultid="8467" heatid="10686" lane="9" entrytime="00:00:32.30" entrycourse="LCM" />
                <RESULT eventid="1373" points="388" swimtime="00:01:10.70" resultid="8468" heatid="10740" lane="8" entrytime="00:01:09.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tayla" lastname="Kalluf Oliveira" birthdate="2011-12-05" gender="F" nation="BRA" license="414583" swrid="5755374" athleteid="8484" externalid="414583">
              <RESULTS>
                <RESULT eventid="1095" points="460" swimtime="00:00:31.63" resultid="8485" heatid="10497" lane="4" entrytime="00:00:33.57" entrycourse="LCM" />
                <RESULT eventid="1147" points="457" swimtime="00:01:07.12" resultid="8486" heatid="10530" lane="2" entrytime="00:01:08.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="437" swimtime="00:00:31.10" resultid="8487" heatid="10606" lane="5" entrytime="00:00:30.81" entrycourse="LCM" />
                <RESULT eventid="1281" points="421" swimtime="00:02:29.65" resultid="8488" heatid="10655" lane="3" entrytime="00:02:38.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                    <SPLIT distance="100" swimtime="00:01:12.43" />
                    <SPLIT distance="150" swimtime="00:01:51.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="384" swimtime="00:01:15.86" resultid="8489" heatid="10701" lane="3" entrytime="00:01:16.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Bulgarelli Castro" birthdate="2012-04-12" gender="M" nation="BRA" license="402125" swrid="5661342" athleteid="8480" externalid="402125">
              <RESULTS>
                <RESULT eventid="1155" points="256" swimtime="00:01:13.06" resultid="8481" heatid="10540" lane="3" entrytime="00:01:12.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="275" swimtime="00:00:32.12" resultid="8482" heatid="10617" lane="8" entrytime="00:00:31.36" entrycourse="LCM" />
                <RESULT eventid="1289" points="266" swimtime="00:02:38.54" resultid="8483" heatid="10662" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                    <SPLIT distance="100" swimtime="00:01:16.29" />
                    <SPLIT distance="150" swimtime="00:01:58.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Bulgarelli Castro" birthdate="2009-04-20" gender="M" nation="BRA" license="401867" swrid="5658058" athleteid="8474" externalid="401867">
              <RESULTS>
                <RESULT eventid="1087" points="283" swimtime="00:03:11.11" resultid="8475" heatid="10488" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.50" />
                    <SPLIT distance="100" swimtime="00:01:29.52" />
                    <SPLIT distance="150" swimtime="00:02:21.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="315" swimtime="00:00:38.13" resultid="8476" heatid="10572" lane="5" entrytime="00:00:38.37" entrycourse="LCM" />
                <RESULT eventid="1155" points="340" swimtime="00:01:06.43" resultid="8477" heatid="10543" lane="6" entrytime="00:01:06.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="330" swimtime="00:00:30.24" resultid="8478" heatid="10620" lane="9" entrytime="00:00:29.74" entrycourse="LCM" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="8479" heatid="10645" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Pascuti Dumke" birthdate="2009-12-28" gender="M" nation="BRA" license="418417" swrid="5706009" athleteid="8495" externalid="418417">
              <RESULTS>
                <RESULT eventid="1155" points="275" swimtime="00:01:11.35" resultid="8496" heatid="10542" lane="2" entrytime="00:01:09.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="303" swimtime="00:00:31.11" resultid="8497" heatid="10617" lane="3" entrytime="00:00:31.02" entrycourse="LCM" />
                <RESULT eventid="1289" points="245" swimtime="00:02:42.99" resultid="8498" heatid="10662" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                    <SPLIT distance="100" swimtime="00:01:15.16" />
                    <SPLIT distance="150" swimtime="00:01:59.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16053" nation="BRA" region="PR" clubid="8546" swrid="93777" name="Fábrica De Nadadores" shortname="Fábrica">
          <ATHLETES>
            <ATHLETE firstname="Gabriel" lastname="Traci Rodrigues" birthdate="2011-03-06" gender="M" nation="BRA" license="406927" swrid="5718893" athleteid="8575" externalid="406927">
              <RESULTS>
                <RESULT eventid="1087" points="202" swimtime="00:03:33.78" resultid="8576" heatid="10487" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.95" />
                    <SPLIT distance="100" swimtime="00:01:39.28" />
                    <SPLIT distance="150" swimtime="00:02:36.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="205" swimtime="00:00:44.01" resultid="8577" heatid="10570" lane="4" entrytime="00:00:45.47" entrycourse="LCM" />
                <RESULT eventid="1155" points="238" swimtime="00:01:14.81" resultid="8578" heatid="10539" lane="2" entrytime="00:01:15.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="252" swimtime="00:00:33.08" resultid="8579" heatid="10614" lane="2" entrytime="00:00:34.06" entrycourse="LCM" />
                <RESULT eventid="1219" points="208" swimtime="00:01:35.98" resultid="8580" heatid="10592" lane="2" entrytime="00:01:41.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="193" swimtime="00:02:56.29" resultid="8581" heatid="10664" lane="6" entrytime="00:03:00.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                    <SPLIT distance="100" swimtime="00:01:16.46" />
                    <SPLIT distance="150" swimtime="00:02:03.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Rumiato Aguilar" birthdate="2011-11-23" gender="M" nation="BRA" license="400277" swrid="5820336" athleteid="8710" externalid="400277">
              <RESULTS>
                <RESULT comment="SW 6.4 - Não começou a executar a virada imediatamente após virar para a posição de peito.  (Horário: 9:41), Na volta dos 50 e 150m." eventid="1071" status="DSQ" swimtime="00:02:47.85" resultid="8711" heatid="10477" lane="0" entrytime="00:02:44.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                    <SPLIT distance="100" swimtime="00:01:19.94" />
                    <SPLIT distance="150" swimtime="00:02:03.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="362" swimtime="00:01:05.09" resultid="8712" heatid="10542" lane="8" entrytime="00:01:09.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="316" swimtime="00:02:29.75" resultid="8713" heatid="10661" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                    <SPLIT distance="100" swimtime="00:01:11.68" />
                    <SPLIT distance="150" swimtime="00:01:50.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="313" swimtime="00:01:15.92" resultid="8714" heatid="10737" lane="2" entrytime="00:01:17.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Magalhães Rezende" birthdate="2010-05-29" gender="F" nation="BRA" license="366960" swrid="5588793" athleteid="8610" externalid="366960">
              <RESULTS>
                <RESULT eventid="1115" points="278" swimtime="00:23:30.09" resultid="8611" heatid="10512" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                    <SPLIT distance="100" swimtime="00:01:19.85" />
                    <SPLIT distance="150" swimtime="00:02:03.69" />
                    <SPLIT distance="200" swimtime="00:02:49.09" />
                    <SPLIT distance="250" swimtime="00:03:35.27" />
                    <SPLIT distance="300" swimtime="00:04:22.10" />
                    <SPLIT distance="350" swimtime="00:05:09.59" />
                    <SPLIT distance="400" swimtime="00:05:57.44" />
                    <SPLIT distance="450" swimtime="00:06:45.35" />
                    <SPLIT distance="500" swimtime="00:07:32.95" />
                    <SPLIT distance="550" swimtime="00:08:20.98" />
                    <SPLIT distance="600" swimtime="00:09:09.24" />
                    <SPLIT distance="650" swimtime="00:09:57.73" />
                    <SPLIT distance="700" swimtime="00:10:45.99" />
                    <SPLIT distance="750" swimtime="00:11:34.11" />
                    <SPLIT distance="800" swimtime="00:12:22.47" />
                    <SPLIT distance="850" swimtime="00:13:11.14" />
                    <SPLIT distance="900" swimtime="00:14:00.12" />
                    <SPLIT distance="950" swimtime="00:14:48.62" />
                    <SPLIT distance="1000" swimtime="00:15:37.63" />
                    <SPLIT distance="1050" swimtime="00:16:26.24" />
                    <SPLIT distance="1100" swimtime="00:17:14.38" />
                    <SPLIT distance="1150" swimtime="00:18:02.90" />
                    <SPLIT distance="1200" swimtime="00:18:49.93" />
                    <SPLIT distance="1250" swimtime="00:19:37.06" />
                    <SPLIT distance="1300" swimtime="00:20:24.07" />
                    <SPLIT distance="1350" swimtime="00:21:11.13" />
                    <SPLIT distance="1400" swimtime="00:21:57.82" />
                    <SPLIT distance="1450" swimtime="00:22:44.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="386" swimtime="00:01:11.01" resultid="8612" heatid="10524" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="268" swimtime="00:12:31.70" resultid="8613" heatid="10633" lane="7" entrytime="00:12:03.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.06" />
                    <SPLIT distance="100" swimtime="00:01:23.91" />
                    <SPLIT distance="150" swimtime="00:02:11.40" />
                    <SPLIT distance="200" swimtime="00:02:59.35" />
                    <SPLIT distance="250" swimtime="00:03:46.97" />
                    <SPLIT distance="300" swimtime="00:04:35.36" />
                    <SPLIT distance="350" swimtime="00:05:22.76" />
                    <SPLIT distance="400" swimtime="00:06:10.47" />
                    <SPLIT distance="450" swimtime="00:06:58.54" />
                    <SPLIT distance="500" swimtime="00:07:46.43" />
                    <SPLIT distance="550" swimtime="00:08:34.71" />
                    <SPLIT distance="600" swimtime="00:09:23.09" />
                    <SPLIT distance="650" swimtime="00:10:10.57" />
                    <SPLIT distance="700" swimtime="00:10:57.88" />
                    <SPLIT distance="750" swimtime="00:11:45.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="402" swimtime="00:00:31.97" resultid="8614" heatid="10600" lane="7" />
                <RESULT eventid="1281" points="353" swimtime="00:02:38.80" resultid="8615" heatid="10653" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                    <SPLIT distance="100" swimtime="00:01:14.29" />
                    <SPLIT distance="150" swimtime="00:01:56.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="314" swimtime="00:05:45.96" resultid="8616" heatid="10712" lane="4" entrytime="00:05:52.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                    <SPLIT distance="100" swimtime="00:01:17.14" />
                    <SPLIT distance="150" swimtime="00:02:00.00" />
                    <SPLIT distance="200" swimtime="00:02:44.32" />
                    <SPLIT distance="250" swimtime="00:03:29.39" />
                    <SPLIT distance="300" swimtime="00:04:15.43" />
                    <SPLIT distance="350" swimtime="00:05:01.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Kenji Yamaguchi" birthdate="2011-08-25" gender="M" nation="BRA" license="385708" swrid="5603862" athleteid="8631" externalid="385708">
              <RESULTS>
                <RESULT eventid="1103" points="361" swimtime="00:00:31.27" resultid="8632" heatid="10503" lane="5" entrytime="00:00:35.21" entrycourse="LCM" />
                <RESULT eventid="1171" points="295" swimtime="00:02:45.70" resultid="8633" heatid="10556" lane="7" entrytime="00:02:54.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.33" />
                    <SPLIT distance="100" swimtime="00:01:16.03" />
                    <SPLIT distance="150" swimtime="00:02:01.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="292" swimtime="00:00:31.50" resultid="8634" heatid="10610" lane="8" />
                <RESULT eventid="1219" points="272" swimtime="00:01:27.71" resultid="8635" heatid="10593" lane="6" entrytime="00:01:30.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="324" swimtime="00:02:45.93" resultid="8636" heatid="10647" lane="1" entrytime="00:02:58.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="100" swimtime="00:01:17.71" />
                    <SPLIT distance="150" swimtime="00:02:07.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="384" swimtime="00:01:08.00" resultid="8637" heatid="10706" lane="3" entrytime="00:01:16.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eloah" lastname="Frasson" birthdate="2012-06-14" gender="F" nation="BRA" license="378338" swrid="5577016" athleteid="8651" externalid="378338">
              <RESULTS>
                <RESULT eventid="1095" points="286" swimtime="00:00:37.06" resultid="8652" heatid="10494" lane="9" />
                <RESULT eventid="1079" points="338" swimtime="00:03:17.37" resultid="8653" heatid="10481" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.77" />
                    <SPLIT distance="100" swimtime="00:01:32.83" />
                    <SPLIT distance="150" swimtime="00:02:26.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="358" swimtime="00:00:41.04" resultid="8654" heatid="10563" lane="0" entrytime="00:00:41.99" entrycourse="LCM" />
                <RESULT eventid="1227" points="323" swimtime="00:00:34.38" resultid="8655" heatid="10602" lane="1" entrytime="00:00:35.66" entrycourse="LCM" />
                <RESULT eventid="1211" points="341" swimtime="00:01:31.71" resultid="8656" heatid="10585" lane="9" entrytime="00:01:34.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="269" swimtime="00:06:04.41" resultid="8657" heatid="10712" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.26" />
                    <SPLIT distance="100" swimtime="00:01:22.42" />
                    <SPLIT distance="150" swimtime="00:02:09.42" />
                    <SPLIT distance="200" swimtime="00:02:56.90" />
                    <SPLIT distance="250" swimtime="00:03:45.27" />
                    <SPLIT distance="300" swimtime="00:04:32.97" />
                    <SPLIT distance="350" swimtime="00:05:20.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rodrigo" lastname="Zanatta Duda" birthdate="2011-09-12" gender="M" nation="BRA" license="406917" swrid="5717307" athleteid="8684" externalid="406917">
              <RESULTS>
                <RESULT eventid="1071" points="377" swimtime="00:02:34.84" resultid="8685" heatid="10477" lane="6" entrytime="00:02:38.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="100" swimtime="00:01:12.29" />
                    <SPLIT distance="150" swimtime="00:01:53.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="210" swimtime="00:00:43.59" resultid="8686" heatid="10571" lane="1" entrytime="00:00:44.11" entrycourse="LCM" />
                <RESULT eventid="1235" points="345" swimtime="00:00:29.81" resultid="8687" heatid="10618" lane="8" entrytime="00:00:30.71" entrycourse="LCM" />
                <RESULT eventid="1305" points="370" swimtime="00:00:32.80" resultid="8688" heatid="10685" lane="5" entrytime="00:00:33.15" entrycourse="LCM" />
                <RESULT eventid="1273" points="300" swimtime="00:02:50.18" resultid="8689" heatid="10647" lane="9" entrytime="00:03:05.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                    <SPLIT distance="100" swimtime="00:01:18.32" />
                    <SPLIT distance="150" swimtime="00:02:10.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="383" swimtime="00:01:11.02" resultid="8690" heatid="10739" lane="5" entrytime="00:01:09.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Moreschi" birthdate="2012-08-09" gender="M" nation="BRA" license="385715" swrid="5603876" athleteid="8617" externalid="385715">
              <RESULTS>
                <RESULT eventid="1103" points="235" swimtime="00:00:36.05" resultid="8618" heatid="10501" lane="8" />
                <RESULT eventid="1187" points="231" swimtime="00:00:42.28" resultid="8619" heatid="10571" lane="8" entrytime="00:00:44.32" entrycourse="LCM" />
                <RESULT eventid="1171" points="180" swimtime="00:03:15.20" resultid="8620" heatid="10555" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.55" />
                    <SPLIT distance="100" swimtime="00:01:35.67" />
                    <SPLIT distance="150" swimtime="00:02:26.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="229" swimtime="00:01:32.96" resultid="8621" heatid="10592" lane="4" entrytime="00:01:38.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="189" swimtime="00:01:26.15" resultid="8622" heatid="10703" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="258" swimtime="00:05:45.42" resultid="8623" heatid="10719" lane="9" entrytime="00:06:25.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                    <SPLIT distance="100" swimtime="00:01:20.31" />
                    <SPLIT distance="150" swimtime="00:02:05.88" />
                    <SPLIT distance="200" swimtime="00:02:51.15" />
                    <SPLIT distance="250" swimtime="00:03:36.49" />
                    <SPLIT distance="300" swimtime="00:04:21.35" />
                    <SPLIT distance="350" swimtime="00:05:05.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jennifer" lastname="De Abreu" birthdate="2009-11-07" gender="F" nation="BRA" license="356212" swrid="5600144" athleteid="8554" externalid="356212">
              <RESULTS>
                <RESULT eventid="1063" points="417" swimtime="00:02:44.74" resultid="8555" heatid="10469" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="340" swimtime="00:02:54.37" resultid="8556" heatid="10554" lane="1" entrytime="00:02:58.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.33" />
                    <SPLIT distance="100" swimtime="00:01:19.98" />
                    <SPLIT distance="150" swimtime="00:02:06.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="489" swimtime="00:00:29.96" resultid="8557" heatid="10608" lane="2" entrytime="00:00:29.54" entrycourse="LCM" />
                <RESULT eventid="1265" points="454" swimtime="00:02:43.99" resultid="8558" heatid="10644" lane="0" entrytime="00:02:42.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.95" />
                    <SPLIT distance="100" swimtime="00:01:19.00" />
                    <SPLIT distance="150" swimtime="00:02:08.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="378" swimtime="00:01:16.30" resultid="8559" heatid="10702" lane="7" entrytime="00:01:12.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="406" swimtime="00:01:17.12" resultid="8560" heatid="10731" lane="6" entrytime="00:01:16.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aline" lastname="Hirano" birthdate="2007-11-13" gender="F" nation="BRA" license="358898" swrid="5622283" athleteid="8677" externalid="358898">
              <RESULTS>
                <RESULT eventid="1115" points="319" swimtime="00:22:25.94" resultid="8678" heatid="10512" lane="3" entrytime="00:20:52.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                    <SPLIT distance="100" swimtime="00:01:19.23" />
                    <SPLIT distance="150" swimtime="00:02:01.99" />
                    <SPLIT distance="200" swimtime="00:02:46.02" />
                    <SPLIT distance="250" swimtime="00:03:29.81" />
                    <SPLIT distance="300" swimtime="00:04:14.94" />
                    <SPLIT distance="350" swimtime="00:05:00.36" />
                    <SPLIT distance="400" swimtime="00:05:46.04" />
                    <SPLIT distance="450" swimtime="00:06:31.75" />
                    <SPLIT distance="500" swimtime="00:07:17.85" />
                    <SPLIT distance="550" swimtime="00:08:01.92" />
                    <SPLIT distance="600" swimtime="00:08:47.02" />
                    <SPLIT distance="650" swimtime="00:09:32.03" />
                    <SPLIT distance="700" swimtime="00:10:17.65" />
                    <SPLIT distance="750" swimtime="00:11:03.02" />
                    <SPLIT distance="800" swimtime="00:11:49.36" />
                    <SPLIT distance="850" swimtime="00:12:35.30" />
                    <SPLIT distance="900" swimtime="00:13:21.17" />
                    <SPLIT distance="950" swimtime="00:14:06.50" />
                    <SPLIT distance="1000" swimtime="00:14:52.70" />
                    <SPLIT distance="1050" swimtime="00:15:37.61" />
                    <SPLIT distance="1100" swimtime="00:16:23.18" />
                    <SPLIT distance="1150" swimtime="00:17:08.43" />
                    <SPLIT distance="1200" swimtime="00:17:53.94" />
                    <SPLIT distance="1250" swimtime="00:18:39.51" />
                    <SPLIT distance="1300" swimtime="00:19:25.91" />
                    <SPLIT distance="1350" swimtime="00:20:12.02" />
                    <SPLIT distance="1400" swimtime="00:20:58.41" />
                    <SPLIT distance="1450" swimtime="00:21:42.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="334" swimtime="00:02:57.34" resultid="8679" heatid="10471" lane="9" entrytime="00:02:56.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.61" />
                    <SPLIT distance="100" swimtime="00:01:24.60" />
                    <SPLIT distance="150" swimtime="00:02:12.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="305" swimtime="00:06:32.76" resultid="8680" heatid="10519" lane="3" entrytime="00:06:08.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.80" />
                    <SPLIT distance="100" swimtime="00:01:38.05" />
                    <SPLIT distance="150" swimtime="00:02:25.77" />
                    <SPLIT distance="200" swimtime="00:03:13.52" />
                    <SPLIT distance="250" swimtime="00:04:13.12" />
                    <SPLIT distance="300" swimtime="00:05:11.26" />
                    <SPLIT distance="350" swimtime="00:05:51.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="324" swimtime="00:11:45.77" resultid="8681" heatid="10632" lane="0" entrytime="00:10:54.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                    <SPLIT distance="100" swimtime="00:01:19.11" />
                    <SPLIT distance="150" swimtime="00:02:01.22" />
                    <SPLIT distance="200" swimtime="00:02:45.39" />
                    <SPLIT distance="250" swimtime="00:03:29.28" />
                    <SPLIT distance="300" swimtime="00:04:14.65" />
                    <SPLIT distance="350" swimtime="00:04:59.44" />
                    <SPLIT distance="400" swimtime="00:05:45.18" />
                    <SPLIT distance="450" swimtime="00:06:29.76" />
                    <SPLIT distance="500" swimtime="00:07:15.56" />
                    <SPLIT distance="550" swimtime="00:08:00.55" />
                    <SPLIT distance="600" swimtime="00:08:46.72" />
                    <SPLIT distance="650" swimtime="00:09:31.82" />
                    <SPLIT distance="700" swimtime="00:10:17.70" />
                    <SPLIT distance="750" swimtime="00:11:01.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="326" swimtime="00:03:03.16" resultid="8682" heatid="10642" lane="8" entrytime="00:02:52.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.52" />
                    <SPLIT distance="100" swimtime="00:01:25.45" />
                    <SPLIT distance="150" swimtime="00:02:22.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="364" swimtime="00:01:19.98" resultid="8683" heatid="10730" lane="5" entrytime="00:01:17.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Arai Junkes" birthdate="2012-08-07" gender="M" nation="BRA" license="424057" athleteid="8741" externalid="424057">
              <RESULTS>
                <RESULT eventid="1103" points="176" swimtime="00:00:39.72" resultid="8742" heatid="10502" lane="0" />
                <RESULT eventid="1155" points="258" swimtime="00:01:12.83" resultid="8743" heatid="10536" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="270" swimtime="00:00:32.33" resultid="8744" heatid="10610" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Zardo" birthdate="2012-05-21" gender="M" nation="BRA" license="423346" swrid="5820329" athleteid="8722" externalid="423346">
              <RESULTS>
                <RESULT eventid="1187" points="142" swimtime="00:00:49.64" resultid="8723" heatid="10570" lane="1" entrytime="00:00:49.76" entrycourse="LCM" />
                <RESULT eventid="1155" points="263" swimtime="00:01:12.37" resultid="8724" heatid="10539" lane="7" entrytime="00:01:15.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="263" swimtime="00:00:32.60" resultid="8725" heatid="10611" lane="1" />
                <RESULT eventid="1219" points="149" swimtime="00:01:47.20" resultid="8726" heatid="10591" lane="4" entrytime="00:01:55.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="253" swimtime="00:02:41.09" resultid="8727" heatid="10664" lane="3" entrytime="00:02:56.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.99" />
                    <SPLIT distance="100" swimtime="00:01:17.65" />
                    <SPLIT distance="150" swimtime="00:02:00.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Pazinato" birthdate="2011-01-05" gender="M" nation="BRA" license="368149" swrid="5603889" athleteid="8638" externalid="368149">
              <RESULTS>
                <RESULT eventid="1071" points="346" swimtime="00:02:39.33" resultid="8639" heatid="10476" lane="2" entrytime="00:02:48.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.03" />
                    <SPLIT distance="100" swimtime="00:01:16.89" />
                    <SPLIT distance="150" swimtime="00:01:57.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="388" swimtime="00:01:03.60" resultid="8640" heatid="10545" lane="4" entrytime="00:01:04.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="398" swimtime="00:00:28.42" resultid="8641" heatid="10619" lane="6" entrytime="00:00:29.85" entrycourse="LCM" />
                <RESULT eventid="1305" points="314" swimtime="00:00:34.62" resultid="8642" heatid="10682" lane="7" />
                <RESULT eventid="1289" points="353" swimtime="00:02:24.19" resultid="8643" heatid="10667" lane="6" entrytime="00:02:29.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.93" />
                    <SPLIT distance="100" swimtime="00:01:07.52" />
                    <SPLIT distance="150" swimtime="00:01:46.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="342" swimtime="00:01:13.75" resultid="8644" heatid="10737" lane="6" entrytime="00:01:16.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucca" lastname="Diedrichs Santos" birthdate="2011-10-27" gender="M" nation="BRA" license="414417" swrid="5755372" athleteid="8698" externalid="414417" />
            <ATHLETE firstname="Luana" lastname="Siqueira Lopes" birthdate="2012-04-28" gender="F" nation="BRA" license="414671" swrid="5755342" athleteid="8735" externalid="414671">
              <RESULTS>
                <RESULT eventid="1095" points="380" swimtime="00:00:33.71" resultid="8736" heatid="10497" lane="2" entrytime="00:00:34.51" entrycourse="LCM" />
                <RESULT eventid="1147" points="410" swimtime="00:01:09.57" resultid="8737" heatid="10529" lane="4" entrytime="00:01:09.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="435" swimtime="00:00:31.15" resultid="8738" heatid="10607" lane="0" entrytime="00:00:30.61" entrycourse="LCM" />
                <RESULT eventid="1281" points="358" swimtime="00:02:38.01" resultid="8739" heatid="10656" lane="0" entrytime="00:02:35.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                    <SPLIT distance="100" swimtime="00:01:14.86" />
                    <SPLIT distance="150" swimtime="00:01:58.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="319" swimtime="00:05:44.43" resultid="8740" heatid="10713" lane="9" entrytime="00:05:51.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.28" />
                    <SPLIT distance="100" swimtime="00:01:20.11" />
                    <SPLIT distance="150" swimtime="00:02:05.56" />
                    <SPLIT distance="200" swimtime="00:02:51.25" />
                    <SPLIT distance="250" swimtime="00:03:35.10" />
                    <SPLIT distance="300" swimtime="00:04:20.48" />
                    <SPLIT distance="350" swimtime="00:05:04.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benicio" lastname="Garcia" birthdate="2011-09-09" gender="M" nation="BRA" license="378347" swrid="5603842" athleteid="8561" externalid="378347">
              <RESULTS>
                <RESULT eventid="1103" points="269" swimtime="00:00:34.46" resultid="8562" heatid="10500" lane="0" />
                <RESULT eventid="1187" points="154" swimtime="00:00:48.40" resultid="8563" heatid="10568" lane="1" />
                <RESULT eventid="1171" points="181" swimtime="00:03:14.98" resultid="8564" heatid="10555" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.75" />
                    <SPLIT distance="100" swimtime="00:01:30.30" />
                    <SPLIT distance="150" swimtime="00:02:21.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="298" swimtime="00:00:31.29" resultid="8565" heatid="10616" lane="9" entrytime="00:00:32.24" entrycourse="LCM" />
                <RESULT eventid="1273" points="225" swimtime="00:03:07.41" resultid="8566" heatid="10646" lane="3" entrytime="00:03:11.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.08" />
                    <SPLIT distance="100" swimtime="00:01:26.35" />
                    <SPLIT distance="150" swimtime="00:02:26.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="217" swimtime="00:01:22.26" resultid="8567" heatid="10705" lane="1" entrytime="00:01:33.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Sales" birthdate="2011-02-28" gender="F" nation="BRA" license="374103" swrid="5616410" athleteid="8645" externalid="374103">
              <RESULTS>
                <RESULT eventid="1095" points="515" swimtime="00:00:30.46" resultid="8646" heatid="10494" lane="2" />
                <RESULT eventid="1163" status="DNS" swimtime="00:00:00.00" resultid="8647" heatid="10553" lane="2" />
                <RESULT eventid="1147" points="484" swimtime="00:01:05.83" resultid="8648" heatid="10531" lane="5" entrytime="00:01:06.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="382" swimtime="00:05:24.18" resultid="8649" heatid="10713" lane="7" entrytime="00:05:37.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                    <SPLIT distance="100" swimtime="00:01:16.40" />
                    <SPLIT distance="150" swimtime="00:01:58.00" />
                    <SPLIT distance="200" swimtime="00:02:39.62" />
                    <SPLIT distance="250" swimtime="00:03:21.49" />
                    <SPLIT distance="300" swimtime="00:04:03.23" />
                    <SPLIT distance="350" swimtime="00:04:44.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="449" swimtime="00:01:12.03" resultid="8650" heatid="10702" lane="1" entrytime="00:01:12.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Britto" birthdate="2012-10-04" gender="M" nation="BRA" license="378350" swrid="5588566" athleteid="8582" externalid="378350">
              <RESULTS>
                <RESULT eventid="1071" points="296" swimtime="00:02:47.82" resultid="8583" heatid="10474" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                    <SPLIT distance="100" swimtime="00:01:21.55" />
                    <SPLIT distance="150" swimtime="00:02:06.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="241" swimtime="00:06:29.16" resultid="8584" heatid="10521" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                    <SPLIT distance="100" swimtime="00:01:28.17" />
                    <SPLIT distance="150" swimtime="00:02:17.80" />
                    <SPLIT distance="200" swimtime="00:03:06.92" />
                    <SPLIT distance="250" swimtime="00:04:02.25" />
                    <SPLIT distance="300" swimtime="00:05:00.23" />
                    <SPLIT distance="350" swimtime="00:05:44.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="319" swimtime="00:00:30.60" resultid="8585" heatid="10614" lane="6" entrytime="00:00:33.67" entrycourse="LCM" />
                <RESULT eventid="1305" points="315" swimtime="00:00:34.61" resultid="8586" heatid="10685" lane="1" entrytime="00:00:35.40" entrycourse="LCM" />
                <RESULT eventid="1273" points="264" swimtime="00:02:57.59" resultid="8587" heatid="10646" lane="2" entrytime="00:03:13.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                    <SPLIT distance="100" swimtime="00:01:22.83" />
                    <SPLIT distance="150" swimtime="00:02:17.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="330" swimtime="00:01:14.65" resultid="8588" heatid="10736" lane="4" entrytime="00:01:20.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Ferreira Rais" birthdate="2007-07-04" gender="M" nation="BRA" license="398656" swrid="5697227" athleteid="8670" externalid="398656">
              <RESULTS>
                <RESULT eventid="1123" points="278" swimtime="00:11:32.35" resultid="8671" heatid="10516" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                    <SPLIT distance="100" swimtime="00:01:11.90" />
                    <SPLIT distance="150" swimtime="00:01:52.94" />
                    <SPLIT distance="200" swimtime="00:02:34.62" />
                    <SPLIT distance="250" swimtime="00:03:18.61" />
                    <SPLIT distance="300" swimtime="00:04:02.23" />
                    <SPLIT distance="350" swimtime="00:04:46.68" />
                    <SPLIT distance="400" swimtime="00:05:31.93" />
                    <SPLIT distance="450" swimtime="00:06:17.15" />
                    <SPLIT distance="500" swimtime="00:07:03.74" />
                    <SPLIT distance="550" swimtime="00:07:49.39" />
                    <SPLIT distance="600" swimtime="00:08:34.68" />
                    <SPLIT distance="650" swimtime="00:09:20.82" />
                    <SPLIT distance="700" swimtime="00:10:06.34" />
                    <SPLIT distance="750" swimtime="00:10:51.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="430" swimtime="00:00:29.50" resultid="8672" heatid="10505" lane="7" entrytime="00:00:31.81" entrycourse="LCM" />
                <RESULT eventid="1155" points="449" swimtime="00:01:00.56" resultid="8673" heatid="10547" lane="6" entrytime="00:01:01.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="465" swimtime="00:00:26.98" resultid="8674" heatid="10623" lane="1" entrytime="00:00:27.68" entrycourse="LCM" />
                <RESULT comment="SW 6.5 - Não terminou a prova enquanto estava de costas.&#10;&#10;&#10;&#10;&#10;&#10;&#10;  (Horário: 16:37), Na volta dos 100m (Costas, Medley Individual)." eventid="1273" status="DSQ" swimtime="00:02:50.58" resultid="8675" heatid="10647" lane="2" entrytime="00:02:57.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="100" swimtime="00:01:17.43" />
                    <SPLIT distance="150" swimtime="00:02:13.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="265" swimtime="00:01:16.92" resultid="8676" heatid="10706" lane="7" entrytime="00:01:17.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="Jose Viana" birthdate="2011-05-25" gender="M" nation="BRA" license="422658" swrid="5820331" athleteid="8705" externalid="422658">
              <RESULTS>
                <RESULT eventid="1187" points="175" swimtime="00:00:46.32" resultid="8706" heatid="10568" lane="5" />
                <RESULT eventid="1155" points="176" swimtime="00:01:22.78" resultid="8707" heatid="10538" lane="3" entrytime="00:01:22.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="189" swimtime="00:00:36.38" resultid="8708" heatid="10613" lane="3" entrytime="00:00:36.57" entrycourse="LCM" />
                <RESULT eventid="1305" points="151" swimtime="00:00:44.13" resultid="8709" heatid="10683" lane="4" entrytime="00:00:43.56" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monique" lastname="Istake" birthdate="2012-04-03" gender="F" nation="BRA" license="372023" swrid="5603857" athleteid="8589" externalid="372023">
              <RESULTS>
                <RESULT eventid="1095" points="394" swimtime="00:00:33.31" resultid="8590" heatid="10497" lane="1" entrytime="00:00:34.94" entrycourse="LCM" />
                <RESULT eventid="1163" points="216" swimtime="00:03:22.92" resultid="8591" heatid="10553" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                    <SPLIT distance="100" swimtime="00:01:29.04" />
                    <SPLIT distance="150" swimtime="00:02:26.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="318" swimtime="00:11:49.72" resultid="8592" heatid="10634" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                    <SPLIT distance="100" swimtime="00:01:16.96" />
                    <SPLIT distance="150" swimtime="00:02:01.42" />
                    <SPLIT distance="200" swimtime="00:02:45.84" />
                    <SPLIT distance="250" swimtime="00:03:30.83" />
                    <SPLIT distance="300" swimtime="00:04:15.32" />
                    <SPLIT distance="350" swimtime="00:05:01.79" />
                    <SPLIT distance="400" swimtime="00:05:48.44" />
                    <SPLIT distance="450" swimtime="00:06:34.67" />
                    <SPLIT distance="500" swimtime="00:07:21.40" />
                    <SPLIT distance="550" swimtime="00:08:06.70" />
                    <SPLIT distance="600" swimtime="00:08:52.41" />
                    <SPLIT distance="650" swimtime="00:09:37.39" />
                    <SPLIT distance="700" swimtime="00:10:23.61" />
                    <SPLIT distance="750" swimtime="00:11:08.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="436" swimtime="00:00:31.12" resultid="8593" heatid="10603" lane="3" entrytime="00:00:33.05" entrycourse="LCM" />
                <RESULT eventid="1281" points="344" swimtime="00:02:40.09" resultid="8594" heatid="10654" lane="4" entrytime="00:02:48.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                    <SPLIT distance="100" swimtime="00:01:15.37" />
                    <SPLIT distance="150" swimtime="00:01:58.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="288" swimtime="00:01:23.54" resultid="8595" heatid="10700" lane="5" entrytime="00:01:26.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruna" lastname="Scalise Drapzichinski" birthdate="2012-03-07" gender="F" nation="BRA" license="378349" swrid="5603909" athleteid="8568" externalid="378349">
              <RESULTS>
                <RESULT eventid="1095" points="392" swimtime="00:00:33.36" resultid="8569" heatid="10496" lane="4" entrytime="00:00:36.49" entrycourse="LCM" />
                <RESULT eventid="1079" points="440" swimtime="00:03:00.82" resultid="8570" heatid="10482" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                    <SPLIT distance="100" swimtime="00:01:23.57" />
                    <SPLIT distance="150" swimtime="00:02:12.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="471" swimtime="00:00:37.47" resultid="8571" heatid="10565" lane="9" entrytime="00:00:37.37" entrycourse="LCM" />
                <RESULT eventid="1147" points="459" swimtime="00:01:07.00" resultid="8572" heatid="10528" lane="4" entrytime="00:01:12.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="465" swimtime="00:00:30.47" resultid="8573" heatid="10606" lane="9" entrytime="00:00:31.19" entrycourse="LCM" />
                <RESULT eventid="1211" points="514" swimtime="00:01:20.02" resultid="8574" heatid="10588" lane="1" entrytime="00:01:22.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Braga" birthdate="2010-05-07" gender="M" nation="BRA" license="378345" swrid="5343953" athleteid="8547" externalid="378345">
              <RESULTS>
                <RESULT eventid="1087" points="481" swimtime="00:02:40.12" resultid="8548" heatid="10491" lane="4" entrytime="00:02:42.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                    <SPLIT distance="100" swimtime="00:01:14.39" />
                    <SPLIT distance="150" swimtime="00:01:57.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="510" swimtime="00:00:32.47" resultid="8549" heatid="10574" lane="2" entrytime="00:00:33.88" entrycourse="LCM" />
                <RESULT eventid="1155" points="369" swimtime="00:01:04.68" resultid="8550" heatid="10544" lane="0" entrytime="00:01:06.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="366" swimtime="00:00:29.22" resultid="8551" heatid="10620" lane="3" entrytime="00:00:29.39" entrycourse="LCM" />
                <RESULT eventid="1219" points="504" swimtime="00:01:11.47" resultid="8552" heatid="10598" lane="8" entrytime="00:01:13.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="398" swimtime="00:02:34.98" resultid="8553" heatid="10648" lane="5" entrytime="00:02:44.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                    <SPLIT distance="100" swimtime="00:01:17.72" />
                    <SPLIT distance="150" swimtime="00:01:58.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benicio" lastname="Alves" birthdate="2012-04-26" gender="M" nation="BRA" license="370588" swrid="5740005" athleteid="8728" externalid="370588">
              <RESULTS>
                <RESULT eventid="1103" status="DNS" swimtime="00:00:00.00" resultid="8729" heatid="10502" lane="2" />
                <RESULT eventid="1155" status="DNS" swimtime="00:00:00.00" resultid="8730" heatid="10538" lane="0" entrytime="00:01:27.75" entrycourse="LCM" />
                <RESULT eventid="1235" status="DNS" swimtime="00:00:00.00" resultid="8731" heatid="10613" lane="6" entrytime="00:00:36.66" entrycourse="LCM" />
                <RESULT eventid="1305" status="DNS" swimtime="00:00:00.00" resultid="8732" heatid="10683" lane="5" entrytime="00:00:44.57" entrycourse="LCM" />
                <RESULT eventid="1289" status="DNS" swimtime="00:00:00.00" resultid="8733" heatid="10664" lane="7" entrytime="00:03:13.01" entrycourse="LCM" />
                <RESULT eventid="1373" status="DNS" swimtime="00:00:00.00" resultid="8734" heatid="10735" lane="3" entrytime="00:01:34.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Rossi" birthdate="2012-05-21" gender="M" nation="BRA" license="378346" swrid="5603901" athleteid="8658" externalid="378346">
              <RESULTS>
                <RESULT eventid="1103" points="205" swimtime="00:00:37.72" resultid="8659" heatid="10502" lane="7" />
                <RESULT eventid="1187" points="170" swimtime="00:00:46.82" resultid="8660" heatid="10566" lane="3" />
                <RESULT eventid="1155" points="277" swimtime="00:01:11.13" resultid="8661" heatid="10540" lane="8" entrytime="00:01:13.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="329" swimtime="00:00:30.26" resultid="8662" heatid="10616" lane="4" entrytime="00:00:31.72" entrycourse="LCM" />
                <RESULT eventid="1305" points="226" swimtime="00:00:38.61" resultid="8663" heatid="10684" lane="3" entrytime="00:00:37.92" entrycourse="LCM" />
                <RESULT eventid="1341" points="174" swimtime="00:01:28.56" resultid="8664" heatid="10704" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="Jacobsen Donati" birthdate="2011-07-14" gender="M" nation="BRA" license="391851" swrid="5615735" athleteid="8624" externalid="391851">
              <RESULTS>
                <RESULT eventid="1071" points="457" swimtime="00:02:25.21" resultid="8625" heatid="10478" lane="8" entrytime="00:02:32.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                    <SPLIT distance="100" swimtime="00:01:09.42" />
                    <SPLIT distance="150" swimtime="00:01:47.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="480" swimtime="00:00:26.69" resultid="8626" heatid="10624" lane="8" entrytime="00:00:27.36" entrycourse="LCM" />
                <RESULT eventid="1305" points="470" swimtime="00:00:30.28" resultid="8627" heatid="10681" lane="1" />
                <RESULT eventid="1289" points="445" swimtime="00:02:13.59" resultid="8628" heatid="10668" lane="1" entrytime="00:02:22.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                    <SPLIT distance="100" swimtime="00:01:04.85" />
                    <SPLIT distance="150" swimtime="00:01:38.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="386" swimtime="00:01:07.91" resultid="8629" heatid="10707" lane="0" entrytime="00:01:15.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="475" swimtime="00:01:06.12" resultid="8630" heatid="10740" lane="2" entrytime="00:01:08.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theodoro" lastname="Marques Serra" birthdate="2009-11-24" gender="M" nation="BRA" license="370661" swrid="5603870" athleteid="8603" externalid="370661">
              <RESULTS>
                <RESULT eventid="1123" points="427" swimtime="00:10:00.28" resultid="8604" heatid="10515" lane="5" entrytime="00:10:20.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                    <SPLIT distance="100" swimtime="00:01:06.23" />
                    <SPLIT distance="150" swimtime="00:01:43.54" />
                    <SPLIT distance="200" swimtime="00:02:21.45" />
                    <SPLIT distance="250" swimtime="00:03:00.12" />
                    <SPLIT distance="300" swimtime="00:03:39.02" />
                    <SPLIT distance="350" swimtime="00:04:17.98" />
                    <SPLIT distance="400" swimtime="00:04:57.03" />
                    <SPLIT distance="450" swimtime="00:05:36.71" />
                    <SPLIT distance="500" swimtime="00:06:15.61" />
                    <SPLIT distance="550" swimtime="00:06:54.08" />
                    <SPLIT distance="600" swimtime="00:07:32.49" />
                    <SPLIT distance="650" swimtime="00:08:10.63" />
                    <SPLIT distance="700" swimtime="00:08:48.64" />
                    <SPLIT distance="750" swimtime="00:09:24.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="405" swimtime="00:00:30.09" resultid="8605" heatid="10499" lane="6" />
                <RESULT eventid="1155" points="458" swimtime="00:01:00.19" resultid="8606" heatid="10546" lane="4" entrytime="00:01:02.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="429" swimtime="00:19:14.25" resultid="8607" heatid="10636" lane="8" entrytime="00:19:29.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                    <SPLIT distance="100" swimtime="00:01:10.74" />
                    <SPLIT distance="150" swimtime="00:01:50.19" />
                    <SPLIT distance="200" swimtime="00:02:28.94" />
                    <SPLIT distance="250" swimtime="00:03:08.61" />
                    <SPLIT distance="300" swimtime="00:03:47.74" />
                    <SPLIT distance="350" swimtime="00:04:27.58" />
                    <SPLIT distance="400" swimtime="00:05:06.76" />
                    <SPLIT distance="450" swimtime="00:05:45.89" />
                    <SPLIT distance="500" swimtime="00:06:24.50" />
                    <SPLIT distance="550" swimtime="00:07:03.85" />
                    <SPLIT distance="600" swimtime="00:07:43.05" />
                    <SPLIT distance="650" swimtime="00:08:22.54" />
                    <SPLIT distance="700" swimtime="00:09:01.51" />
                    <SPLIT distance="750" swimtime="00:09:40.83" />
                    <SPLIT distance="800" swimtime="00:10:19.76" />
                    <SPLIT distance="850" swimtime="00:10:58.56" />
                    <SPLIT distance="900" swimtime="00:11:36.93" />
                    <SPLIT distance="950" swimtime="00:12:16.45" />
                    <SPLIT distance="1000" swimtime="00:12:54.80" />
                    <SPLIT distance="1050" swimtime="00:13:33.85" />
                    <SPLIT distance="1100" swimtime="00:14:12.30" />
                    <SPLIT distance="1150" swimtime="00:14:51.30" />
                    <SPLIT distance="1200" swimtime="00:15:29.28" />
                    <SPLIT distance="1250" swimtime="00:16:07.68" />
                    <SPLIT distance="1300" swimtime="00:16:45.48" />
                    <SPLIT distance="1350" swimtime="00:17:23.24" />
                    <SPLIT distance="1400" swimtime="00:18:00.86" />
                    <SPLIT distance="1450" swimtime="00:18:38.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="453" swimtime="00:02:12.81" resultid="8608" heatid="10670" lane="1" entrytime="00:02:17.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.05" />
                    <SPLIT distance="100" swimtime="00:01:02.07" />
                    <SPLIT distance="150" swimtime="00:01:37.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="410" swimtime="00:01:09.45" resultid="8609" heatid="10740" lane="9" entrytime="00:01:09.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernanda" lastname="Camillo Sabim" birthdate="2010-08-02" gender="F" nation="BRA" license="406931" swrid="5723021" athleteid="8691" externalid="406931">
              <RESULTS>
                <RESULT eventid="1079" points="369" swimtime="00:03:11.61" resultid="8692" heatid="10483" lane="8" entrytime="00:03:17.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                    <SPLIT distance="100" swimtime="00:01:30.82" />
                    <SPLIT distance="150" swimtime="00:02:21.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="345" swimtime="00:00:41.56" resultid="8693" heatid="10563" lane="1" entrytime="00:00:41.57" entrycourse="LCM" />
                <RESULT eventid="1147" points="369" swimtime="00:01:12.08" resultid="8694" heatid="10528" lane="6" entrytime="00:01:12.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="359" swimtime="00:01:30.20" resultid="8695" heatid="10585" lane="4" entrytime="00:01:31.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="319" swimtime="00:00:39.29" resultid="8696" heatid="10678" lane="2" entrytime="00:00:41.20" entrycourse="LCM" />
                <RESULT eventid="1365" points="322" swimtime="00:01:23.31" resultid="8697" heatid="10728" lane="7" entrytime="00:01:27.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Ribeiro Melo" birthdate="2011-07-01" gender="F" nation="BRA" license="390923" swrid="5602577" athleteid="8596" externalid="390923">
              <RESULTS>
                <RESULT eventid="1179" points="303" swimtime="00:00:43.38" resultid="8597" heatid="10562" lane="3" entrytime="00:00:43.97" entrycourse="LCM" />
                <RESULT eventid="1147" points="450" swimtime="00:01:07.44" resultid="8598" heatid="10531" lane="6" entrytime="00:01:07.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="474" swimtime="00:00:30.26" resultid="8599" heatid="10607" lane="2" entrytime="00:00:30.25" entrycourse="LCM" />
                <RESULT eventid="1281" points="370" swimtime="00:02:36.28" resultid="8600" heatid="10658" lane="3" entrytime="00:02:24.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                    <SPLIT distance="100" swimtime="00:01:13.59" />
                    <SPLIT distance="150" swimtime="00:01:55.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="412" swimtime="00:05:16.22" resultid="8601" heatid="10714" lane="0" entrytime="00:05:28.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                    <SPLIT distance="100" swimtime="00:01:12.99" />
                    <SPLIT distance="150" swimtime="00:01:52.93" />
                    <SPLIT distance="200" swimtime="00:02:34.23" />
                    <SPLIT distance="250" swimtime="00:03:15.39" />
                    <SPLIT distance="300" swimtime="00:03:56.76" />
                    <SPLIT distance="350" swimtime="00:04:37.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="345" swimtime="00:01:21.38" resultid="8602" heatid="10729" lane="7" entrytime="00:01:24.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emanuele" lastname="De Vieira" birthdate="2011-02-04" gender="F" nation="BRA" license="422791" swrid="5820334" athleteid="8715" externalid="422791">
              <RESULTS>
                <RESULT eventid="1095" points="186" swimtime="00:00:42.75" resultid="8716" heatid="10495" lane="4" entrytime="00:00:44.23" entrycourse="LCM" />
                <RESULT eventid="1179" points="226" swimtime="00:00:47.82" resultid="8717" heatid="10561" lane="9" />
                <RESULT eventid="1147" points="289" swimtime="00:01:18.18" resultid="8718" heatid="10526" lane="0" entrytime="00:01:20.88" entrycourse="LCM" />
                <RESULT eventid="1227" points="211" swimtime="00:00:39.65" resultid="8719" heatid="10600" lane="4" />
                <RESULT eventid="1297" points="206" swimtime="00:00:45.41" resultid="8720" heatid="10676" lane="6" />
                <RESULT eventid="1365" points="196" swimtime="00:01:38.29" resultid="8721" heatid="10727" lane="9" entrytime="00:01:38.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Livia" lastname="Eloisa Silva" birthdate="2012-03-03" gender="F" nation="BRA" license="399725" swrid="5651341" athleteid="8665" externalid="399725">
              <RESULTS>
                <RESULT eventid="1147" points="185" swimtime="00:01:30.72" resultid="8666" heatid="10525" lane="0" />
                <RESULT eventid="1227" points="181" swimtime="00:00:41.67" resultid="8667" heatid="10601" lane="1" />
                <RESULT eventid="1297" points="228" swimtime="00:00:43.91" resultid="8668" heatid="10677" lane="3" />
                <RESULT eventid="1365" points="205" swimtime="00:01:36.81" resultid="8669" heatid="10726" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ian" lastname="Thierbach Ruiz" birthdate="2011-10-12" gender="M" nation="BRA" license="413946" swrid="5755380" athleteid="8699" externalid="413946">
              <RESULTS>
                <RESULT eventid="1103" points="257" swimtime="00:00:35.00" resultid="8700" heatid="10503" lane="2" entrytime="00:00:35.90" entrycourse="LCM" />
                <RESULT eventid="1187" points="260" swimtime="00:00:40.61" resultid="8701" heatid="10570" lane="2" entrytime="00:00:47.86" entrycourse="LCM" />
                <RESULT eventid="1235" points="287" swimtime="00:00:31.67" resultid="8702" heatid="10615" lane="0" entrytime="00:00:33.25" entrycourse="LCM" />
                <RESULT eventid="1273" points="265" swimtime="00:02:57.46" resultid="8703" heatid="10645" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="100" swimtime="00:01:21.26" />
                    <SPLIT distance="150" swimtime="00:02:17.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="186" swimtime="00:01:26.58" resultid="8704" heatid="10705" lane="3" entrytime="00:01:25.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="14" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1203" points="331" swimtime="00:10:04.97" resultid="8749" heatid="10579" lane="6" entrytime="00:10:32.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.25" />
                    <SPLIT distance="100" swimtime="00:01:02.56" />
                    <SPLIT distance="150" swimtime="00:01:38.62" />
                    <SPLIT distance="200" swimtime="00:02:15.10" />
                    <SPLIT distance="250" swimtime="00:02:48.80" />
                    <SPLIT distance="300" swimtime="00:03:30.94" />
                    <SPLIT distance="350" swimtime="00:04:13.85" />
                    <SPLIT distance="400" swimtime="00:04:54.98" />
                    <SPLIT distance="450" swimtime="00:05:27.58" />
                    <SPLIT distance="500" swimtime="00:06:09.31" />
                    <SPLIT distance="550" swimtime="00:06:55.01" />
                    <SPLIT distance="600" swimtime="00:07:37.84" />
                    <SPLIT distance="700" swimtime="00:08:44.10" />
                    <SPLIT distance="750" swimtime="00:09:24.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8624" number="1" />
                    <RELAYPOSITION athleteid="8684" number="2" />
                    <RELAYPOSITION athleteid="8582" number="3" />
                    <RELAYPOSITION athleteid="8638" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1323" points="252" swimtime="00:05:27.31" resultid="8750" heatid="10693" lane="2" entrytime="00:05:47.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                    <SPLIT distance="100" swimtime="00:01:15.99" />
                    <SPLIT distance="150" swimtime="00:01:58.26" />
                    <SPLIT distance="200" swimtime="00:02:47.08" />
                    <SPLIT distance="250" swimtime="00:03:25.45" />
                    <SPLIT distance="300" swimtime="00:04:15.46" />
                    <SPLIT distance="350" swimtime="00:04:49.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8582" number="1" />
                    <RELAYPOSITION athleteid="8617" number="2" />
                    <RELAYPOSITION athleteid="8658" number="3" />
                    <RELAYPOSITION athleteid="8722" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1391" points="292" swimtime="00:04:43.51" resultid="8753" heatid="10748" lane="1" entrytime="00:05:02.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.64" />
                    <SPLIT distance="100" swimtime="00:01:13.03" />
                    <SPLIT distance="150" swimtime="00:01:46.65" />
                    <SPLIT distance="200" swimtime="00:02:26.55" />
                    <SPLIT distance="250" swimtime="00:02:58.04" />
                    <SPLIT distance="300" swimtime="00:03:35.22" />
                    <SPLIT distance="350" swimtime="00:04:07.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8722" number="1" />
                    <RELAYPOSITION athleteid="8617" number="2" />
                    <RELAYPOSITION athleteid="8582" number="3" />
                    <RELAYPOSITION athleteid="8658" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1325" points="358" swimtime="00:04:51.06" resultid="8751" heatid="10695" lane="1" entrytime="00:05:47.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                    <SPLIT distance="100" swimtime="00:01:11.97" />
                    <SPLIT distance="150" swimtime="00:01:53.44" />
                    <SPLIT distance="200" swimtime="00:02:39.58" />
                    <SPLIT distance="250" swimtime="00:03:11.87" />
                    <SPLIT distance="300" swimtime="00:03:49.89" />
                    <SPLIT distance="350" swimtime="00:04:17.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8684" number="1" />
                    <RELAYPOSITION athleteid="8631" number="2" />
                    <RELAYPOSITION athleteid="8624" number="3" />
                    <RELAYPOSITION athleteid="8638" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1393" points="391" swimtime="00:04:17.33" resultid="8752" heatid="10750" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.25" />
                    <SPLIT distance="100" swimtime="00:00:58.81" />
                    <SPLIT distance="150" swimtime="00:01:29.46" />
                    <SPLIT distance="200" swimtime="00:02:05.04" />
                    <SPLIT distance="250" swimtime="00:02:36.53" />
                    <SPLIT distance="300" swimtime="00:03:13.87" />
                    <SPLIT distance="350" swimtime="00:03:43.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8624" number="1" />
                    <RELAYPOSITION athleteid="8710" number="2" />
                    <RELAYPOSITION athleteid="8684" number="3" />
                    <RELAYPOSITION athleteid="8638" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="FÁBRICA DE NADADORES &quot;B&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1325" status="DNS" swimtime="00:00:00.00" resultid="8757" heatid="10695" lane="8">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8710" number="1" />
                    <RELAYPOSITION athleteid="8699" number="2" />
                    <RELAYPOSITION athleteid="8561" number="3" />
                    <RELAYPOSITION athleteid="8575" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1393" points="283" swimtime="00:04:46.69" resultid="8758" heatid="10749" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                    <SPLIT distance="100" swimtime="00:01:11.80" />
                    <SPLIT distance="150" swimtime="00:01:46.49" />
                    <SPLIT distance="200" swimtime="00:02:25.23" />
                    <SPLIT distance="250" swimtime="00:02:57.18" />
                    <SPLIT distance="300" swimtime="00:03:35.23" />
                    <SPLIT distance="350" swimtime="00:04:08.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8561" number="1" />
                    <RELAYPOSITION athleteid="8575" number="2" />
                    <RELAYPOSITION athleteid="8699" number="3" />
                    <RELAYPOSITION athleteid="8631" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1195" points="371" swimtime="00:10:36.34" resultid="8745" heatid="10576" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.62" />
                    <SPLIT distance="100" swimtime="00:01:15.20" />
                    <SPLIT distance="150" swimtime="00:01:56.58" />
                    <SPLIT distance="200" swimtime="00:02:34.12" />
                    <SPLIT distance="250" swimtime="00:03:07.58" />
                    <SPLIT distance="300" swimtime="00:03:48.28" />
                    <SPLIT distance="350" swimtime="00:04:30.63" />
                    <SPLIT distance="400" swimtime="00:05:13.91" />
                    <SPLIT distance="450" swimtime="00:05:50.71" />
                    <SPLIT distance="500" swimtime="00:06:34.90" />
                    <SPLIT distance="550" swimtime="00:07:19.89" />
                    <SPLIT distance="600" swimtime="00:07:59.09" />
                    <SPLIT distance="650" swimtime="00:08:36.01" />
                    <SPLIT distance="700" swimtime="00:09:17.83" />
                    <SPLIT distance="750" swimtime="00:09:59.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8596" number="1" />
                    <RELAYPOSITION athleteid="8568" number="2" />
                    <RELAYPOSITION athleteid="8589" number="3" />
                    <RELAYPOSITION athleteid="8735" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1313" points="363" swimtime="00:05:21.84" resultid="8746" heatid="10688" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                    <SPLIT distance="100" swimtime="00:01:19.38" />
                    <SPLIT distance="150" swimtime="00:01:59.55" />
                    <SPLIT distance="200" swimtime="00:02:48.02" />
                    <SPLIT distance="250" swimtime="00:03:24.54" />
                    <SPLIT distance="350" swimtime="00:04:43.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8568" number="1" />
                    <RELAYPOSITION athleteid="8651" number="2" />
                    <RELAYPOSITION athleteid="8589" number="3" />
                    <RELAYPOSITION athleteid="8735" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1381" points="394" swimtime="00:04:43.67" resultid="8747" heatid="10743" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                    <SPLIT distance="100" swimtime="00:01:10.22" />
                    <SPLIT distance="150" swimtime="00:01:45.20" />
                    <SPLIT distance="200" swimtime="00:02:25.03" />
                    <SPLIT distance="250" swimtime="00:02:55.96" />
                    <SPLIT distance="300" swimtime="00:03:32.86" />
                    <SPLIT distance="350" swimtime="00:04:04.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8735" number="1" />
                    <RELAYPOSITION athleteid="8651" number="2" />
                    <RELAYPOSITION athleteid="8568" number="3" />
                    <RELAYPOSITION athleteid="8589" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1383" points="321" swimtime="00:05:03.71" resultid="8748" heatid="10744" lane="7" entrytime="00:05:07.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:01:08.72" />
                    <SPLIT distance="150" swimtime="00:01:44.21" />
                    <SPLIT distance="200" swimtime="00:02:25.90" />
                    <SPLIT distance="250" swimtime="00:03:08.92" />
                    <SPLIT distance="300" swimtime="00:03:58.07" />
                    <SPLIT distance="350" swimtime="00:04:28.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8596" number="1" />
                    <RELAYPOSITION athleteid="8715" number="2" />
                    <RELAYPOSITION athleteid="8665" number="3" />
                    <RELAYPOSITION athleteid="8645" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1113" points="401" swimtime="00:04:54.79" resultid="8754" heatid="10510" lane="1" entrytime="00:05:45.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                    <SPLIT distance="150" swimtime="00:01:46.70" />
                    <SPLIT distance="250" swimtime="00:03:06.39" />
                    <SPLIT distance="300" swimtime="00:03:47.09" />
                    <SPLIT distance="350" swimtime="00:04:18.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8624" number="1" />
                    <RELAYPOSITION athleteid="8631" number="2" />
                    <RELAYPOSITION athleteid="8645" number="3" />
                    <RELAYPOSITION athleteid="8596" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="X" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1111" points="346" swimtime="00:05:09.42" resultid="8755" heatid="10509" lane="2" entrytime="00:05:29.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                    <SPLIT distance="100" swimtime="00:01:14.86" />
                    <SPLIT distance="150" swimtime="00:01:51.29" />
                    <SPLIT distance="200" swimtime="00:02:37.07" />
                    <SPLIT distance="250" swimtime="00:03:13.06" />
                    <SPLIT distance="300" swimtime="00:04:00.25" />
                    <SPLIT distance="350" swimtime="00:04:32.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8582" number="1" />
                    <RELAYPOSITION athleteid="8568" number="2" />
                    <RELAYPOSITION athleteid="8589" number="3" />
                    <RELAYPOSITION athleteid="8658" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="X" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1245" points="453" swimtime="00:04:42.97" resultid="8756" heatid="10630" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                    <SPLIT distance="100" swimtime="00:01:09.17" />
                    <SPLIT distance="150" swimtime="00:01:42.35" />
                    <SPLIT distance="200" swimtime="00:02:21.07" />
                    <SPLIT distance="250" swimtime="00:02:54.06" />
                    <SPLIT distance="300" swimtime="00:03:34.23" />
                    <SPLIT distance="350" swimtime="00:04:06.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8603" number="1" />
                    <RELAYPOSITION athleteid="8547" number="2" />
                    <RELAYPOSITION athleteid="8554" number="3" />
                    <RELAYPOSITION athleteid="8610" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="X" name="FÁBRICA DE NADADORES &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1111" points="262" swimtime="00:05:39.78" resultid="8759" heatid="10509" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.60" />
                    <SPLIT distance="100" swimtime="00:01:33.35" />
                    <SPLIT distance="150" swimtime="00:02:14.17" />
                    <SPLIT distance="200" swimtime="00:03:03.47" />
                    <SPLIT distance="250" swimtime="00:03:39.93" />
                    <SPLIT distance="300" swimtime="00:04:28.68" />
                    <SPLIT distance="350" swimtime="00:05:02.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8735" number="1" />
                    <RELAYPOSITION athleteid="8651" number="2" />
                    <RELAYPOSITION athleteid="8617" number="3" />
                    <RELAYPOSITION athleteid="8722" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="19586" nation="BRA" region="PR" clubid="9495" swrid="95625" name="Winners Vanguarda Gestao Esportiva E Competitiva" shortname="Winners">
          <ATHLETES>
            <ATHLETE firstname="Guilherme" lastname="Kerniski Demantova" birthdate="1982-05-25" gender="M" nation="BRA" license="398222" swrid="5653293" athleteid="9555" externalid="398222" level="DKMBANK">
              <RESULTS>
                <RESULT eventid="1123" points="398" swimtime="00:10:14.63" resultid="9556" heatid="10515" lane="3" entrytime="00:10:20.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                    <SPLIT distance="100" swimtime="00:01:12.54" />
                    <SPLIT distance="150" swimtime="00:01:50.79" />
                    <SPLIT distance="200" swimtime="00:02:29.42" />
                    <SPLIT distance="250" swimtime="00:03:08.12" />
                    <SPLIT distance="300" swimtime="00:03:46.82" />
                    <SPLIT distance="350" swimtime="00:04:25.46" />
                    <SPLIT distance="400" swimtime="00:05:04.46" />
                    <SPLIT distance="450" swimtime="00:05:43.29" />
                    <SPLIT distance="500" swimtime="00:06:22.58" />
                    <SPLIT distance="550" swimtime="00:07:01.47" />
                    <SPLIT distance="600" swimtime="00:07:40.57" />
                    <SPLIT distance="650" swimtime="00:08:19.41" />
                    <SPLIT distance="700" swimtime="00:08:58.72" />
                    <SPLIT distance="750" swimtime="00:09:37.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="301" swimtime="00:06:01.61" resultid="9557" heatid="10521" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.81" />
                    <SPLIT distance="100" swimtime="00:01:26.77" />
                    <SPLIT distance="200" swimtime="00:03:06.73" />
                    <SPLIT distance="250" swimtime="00:03:57.42" />
                    <SPLIT distance="300" swimtime="00:04:46.87" />
                    <SPLIT distance="350" swimtime="00:05:25.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="361" swimtime="00:20:22.38" resultid="9558" heatid="10637" lane="3" entrytime="00:20:14.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.14" />
                    <SPLIT distance="100" swimtime="00:01:20.74" />
                    <SPLIT distance="150" swimtime="00:02:02.60" />
                    <SPLIT distance="200" swimtime="00:02:45.39" />
                    <SPLIT distance="250" swimtime="00:03:27.28" />
                    <SPLIT distance="300" swimtime="00:04:10.21" />
                    <SPLIT distance="350" swimtime="00:04:51.82" />
                    <SPLIT distance="400" swimtime="00:05:33.66" />
                    <SPLIT distance="450" swimtime="00:06:14.88" />
                    <SPLIT distance="500" swimtime="00:06:56.87" />
                    <SPLIT distance="550" swimtime="00:07:37.80" />
                    <SPLIT distance="600" swimtime="00:08:19.47" />
                    <SPLIT distance="650" swimtime="00:09:00.74" />
                    <SPLIT distance="700" swimtime="00:09:42.59" />
                    <SPLIT distance="750" swimtime="00:10:23.24" />
                    <SPLIT distance="800" swimtime="00:11:04.87" />
                    <SPLIT distance="850" swimtime="00:11:45.60" />
                    <SPLIT distance="900" swimtime="00:12:26.74" />
                    <SPLIT distance="950" swimtime="00:13:06.71" />
                    <SPLIT distance="1000" swimtime="00:13:47.88" />
                    <SPLIT distance="1050" swimtime="00:14:28.08" />
                    <SPLIT distance="1100" swimtime="00:15:08.43" />
                    <SPLIT distance="1150" swimtime="00:15:48.19" />
                    <SPLIT distance="1200" swimtime="00:16:28.21" />
                    <SPLIT distance="1250" swimtime="00:17:07.69" />
                    <SPLIT distance="1300" swimtime="00:17:47.45" />
                    <SPLIT distance="1350" swimtime="00:18:26.79" />
                    <SPLIT distance="1400" swimtime="00:19:06.10" />
                    <SPLIT distance="1450" swimtime="00:19:44.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="417" swimtime="00:02:16.45" resultid="9559" heatid="10668" lane="5" entrytime="00:02:21.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.82" />
                    <SPLIT distance="100" swimtime="00:01:05.94" />
                    <SPLIT distance="150" swimtime="00:01:41.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="424" swimtime="00:04:52.79" resultid="9560" heatid="10720" lane="4" entrytime="00:04:59.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                    <SPLIT distance="100" swimtime="00:01:08.77" />
                    <SPLIT distance="150" swimtime="00:01:45.66" />
                    <SPLIT distance="200" swimtime="00:02:22.92" />
                    <SPLIT distance="250" swimtime="00:03:00.24" />
                    <SPLIT distance="300" swimtime="00:03:38.16" />
                    <SPLIT distance="350" swimtime="00:04:16.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="211" swimtime="00:01:26.58" resultid="9561" heatid="10733" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karine" lastname="Correa" birthdate="2002-08-01" gender="F" nation="BRA" license="385191" swrid="5600141" athleteid="9574" externalid="385191">
              <RESULTS>
                <RESULT eventid="1095" points="267" swimtime="00:00:37.91" resultid="9575" heatid="10495" lane="1" />
                <RESULT eventid="1147" points="367" swimtime="00:01:12.20" resultid="9576" heatid="10529" lane="0" entrytime="00:01:12.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="244" swimtime="00:12:54.99" resultid="9577" heatid="10633" lane="1" entrytime="00:12:19.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.56" />
                    <SPLIT distance="100" swimtime="00:01:22.90" />
                    <SPLIT distance="150" swimtime="00:02:10.03" />
                    <SPLIT distance="200" swimtime="00:02:58.56" />
                    <SPLIT distance="250" swimtime="00:03:47.16" />
                    <SPLIT distance="300" swimtime="00:04:37.17" />
                    <SPLIT distance="350" swimtime="00:05:27.16" />
                    <SPLIT distance="400" swimtime="00:06:18.34" />
                    <SPLIT distance="450" swimtime="00:07:09.44" />
                    <SPLIT distance="500" swimtime="00:07:59.95" />
                    <SPLIT distance="550" swimtime="00:08:49.88" />
                    <SPLIT distance="600" swimtime="00:09:39.81" />
                    <SPLIT distance="650" swimtime="00:10:29.50" />
                    <SPLIT distance="700" swimtime="00:11:19.48" />
                    <SPLIT distance="750" swimtime="00:12:08.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="374" swimtime="00:00:32.76" resultid="9578" heatid="10604" lane="7" entrytime="00:00:32.22" entrycourse="LCM" />
                <RESULT eventid="1281" points="325" swimtime="00:02:43.19" resultid="9579" heatid="10655" lane="7" entrytime="00:02:42.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.48" />
                    <SPLIT distance="100" swimtime="00:01:17.62" />
                    <SPLIT distance="150" swimtime="00:02:01.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="275" swimtime="00:06:01.81" resultid="9580" heatid="10713" lane="1" entrytime="00:05:42.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.15" />
                    <SPLIT distance="100" swimtime="00:01:18.99" />
                    <SPLIT distance="150" swimtime="00:02:02.87" />
                    <SPLIT distance="200" swimtime="00:02:49.40" />
                    <SPLIT distance="250" swimtime="00:03:37.14" />
                    <SPLIT distance="300" swimtime="00:04:25.81" />
                    <SPLIT distance="350" swimtime="00:05:14.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose" lastname="Salazar" birthdate="1989-06-25" gender="M" nation="BRA" license="99446" swrid="5811238" athleteid="9597" externalid="99446" level="DKMBANK">
              <RESULTS>
                <RESULT eventid="1103" points="310" swimtime="00:00:32.88" resultid="9598" heatid="10501" lane="5" />
                <RESULT eventid="1087" points="248" swimtime="00:03:19.48" resultid="9599" heatid="10488" lane="6" entrytime="00:03:26.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.19" />
                    <SPLIT distance="100" swimtime="00:01:38.32" />
                    <SPLIT distance="150" swimtime="00:02:32.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="346" swimtime="00:00:36.95" resultid="9600" heatid="10573" lane="9" entrytime="00:00:36.92" entrycourse="LCM" />
                <RESULT eventid="1219" points="291" swimtime="00:01:25.76" resultid="9601" heatid="10593" lane="5" entrytime="00:01:29.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.88" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.4 - Movimentos das pernas não simultâneos.  (Horário: 16:27), Peito, Medley Individual." eventid="1273" status="DSQ" swimtime="00:02:57.39" resultid="9602" heatid="10645" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                    <SPLIT distance="100" swimtime="00:01:21.15" />
                    <SPLIT distance="150" swimtime="00:02:15.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Araujo" birthdate="2003-11-09" gender="M" nation="BRA" license="307551" swrid="5820327" athleteid="9543" externalid="307551" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1103" points="492" swimtime="00:00:28.20" resultid="9544" heatid="10507" lane="4" entrytime="00:00:27.70" entrycourse="LCM" />
                <RESULT eventid="1155" points="593" swimtime="00:00:55.21" resultid="9545" heatid="10551" lane="5" entrytime="00:00:55.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="546" swimtime="00:00:25.57" resultid="9546" heatid="10627" lane="1" entrytime="00:00:25.25" entrycourse="LCM" />
                <RESULT eventid="1289" points="506" swimtime="00:02:07.99" resultid="9547" heatid="10663" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.56" />
                    <SPLIT distance="100" swimtime="00:01:01.54" />
                    <SPLIT distance="150" swimtime="00:01:35.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="480" swimtime="00:01:03.13" resultid="9548" heatid="10704" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Zanatta Flizikowski" birthdate="2010-01-08" gender="F" nation="BRA" license="367051" swrid="5588969" athleteid="9585" externalid="367051">
              <RESULTS>
                <RESULT eventid="1095" points="331" swimtime="00:00:35.31" resultid="9586" heatid="10497" lane="3" entrytime="00:00:34.27" entrycourse="LCM" />
                <RESULT eventid="1147" points="411" swimtime="00:01:09.50" resultid="9587" heatid="10531" lane="4" entrytime="00:01:06.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="416" swimtime="00:00:31.62" resultid="9588" heatid="10605" lane="1" entrytime="00:00:31.43" entrycourse="LCM" />
                <RESULT comment="SW 10.2 - Não completou a distância total da prova.  (Horário: 17:15)" eventid="1281" status="DSQ" swimtime="00:00:00.00" resultid="9589" heatid="10656" lane="3" entrytime="00:02:32.14" entrycourse="LCM" />
                <RESULT eventid="1333" points="241" swimtime="00:01:28.65" resultid="9590" heatid="10701" lane="9" entrytime="00:01:23.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Carvalho Rodrigues" birthdate="2004-01-17" gender="F" nation="BRA" license="249307" swrid="5820338" athleteid="9524" externalid="249307">
              <RESULTS>
                <RESULT eventid="1179" points="389" swimtime="00:00:39.93" resultid="9525" heatid="10563" lane="5" entrytime="00:00:40.76" entrycourse="LCM" />
                <RESULT eventid="1147" points="397" swimtime="00:01:10.30" resultid="9526" heatid="10528" lane="5" entrytime="00:01:12.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="436" swimtime="00:00:31.13" resultid="9527" heatid="10606" lane="7" entrytime="00:00:30.97" entrycourse="LCM" />
                <RESULT eventid="1211" points="335" swimtime="00:01:32.29" resultid="9528" heatid="10583" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="299" swimtime="00:00:40.15" resultid="9529" heatid="10675" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mauricio" lastname="Furtado Niwa" birthdate="1978-05-30" gender="M" nation="BRA" license="398757" swrid="5653291" athleteid="9569" externalid="398757" level="DKMBANK">
              <RESULTS>
                <RESULT eventid="1171" points="343" swimtime="00:02:37.62" resultid="9570" heatid="10557" lane="3" entrytime="00:02:31.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                    <SPLIT distance="100" swimtime="00:01:15.18" />
                    <SPLIT distance="150" swimtime="00:01:57.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="498" swimtime="00:00:26.37" resultid="9571" heatid="10625" lane="8" entrytime="00:00:26.83" entrycourse="LCM" />
                <RESULT eventid="1289" points="447" swimtime="00:02:13.37" resultid="9572" heatid="10671" lane="6" entrytime="00:02:11.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.08" />
                    <SPLIT distance="100" swimtime="00:01:04.63" />
                    <SPLIT distance="150" swimtime="00:01:39.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="504" swimtime="00:01:02.13" resultid="9573" heatid="10710" lane="6" entrytime="00:01:02.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="De Almeida Figueiredo" birthdate="1998-08-25" gender="M" nation="BRA" license="151442" swrid="5820339" athleteid="9496" externalid="151442">
              <RESULTS>
                <RESULT eventid="1155" points="563" swimtime="00:00:56.17" resultid="9497" heatid="10550" lane="3" entrytime="00:00:56.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="535" swimtime="00:00:25.75" resultid="9498" heatid="10626" lane="8" entrytime="00:00:25.96" entrycourse="LCM" />
                <RESULT eventid="1373" points="418" swimtime="00:01:08.99" resultid="9499" heatid="10733" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Allana" lastname="Lacerda" birthdate="2005-03-15" gender="F" nation="BRA" license="295186" swrid="5600197" athleteid="9530" externalid="295186" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1079" points="414" swimtime="00:03:04.44" resultid="9531" heatid="10485" lane="0" entrytime="00:03:02.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.57" />
                    <SPLIT distance="100" swimtime="00:01:28.59" />
                    <SPLIT distance="150" swimtime="00:02:15.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="423" swimtime="00:00:38.84" resultid="9532" heatid="10564" lane="7" entrytime="00:00:38.84" entrycourse="LCM" />
                <RESULT eventid="1211" points="403" swimtime="00:01:26.78" resultid="9533" heatid="10587" lane="5" entrytime="00:01:24.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.49" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.4 - Movimentos das pernas não simultâneos.  (Horário: 16:18),  Peito, Medley Individual." eventid="1265" status="DSQ" swimtime="00:02:48.35" resultid="9534" heatid="10643" lane="8" entrytime="00:02:46.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                    <SPLIT distance="100" swimtime="00:01:21.80" />
                    <SPLIT distance="150" swimtime="00:02:08.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="373" swimtime="00:05:26.74" resultid="9535" heatid="10714" lane="7" entrytime="00:05:18.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                    <SPLIT distance="100" swimtime="00:01:17.63" />
                    <SPLIT distance="150" swimtime="00:01:59.62" />
                    <SPLIT distance="200" swimtime="00:02:41.80" />
                    <SPLIT distance="250" swimtime="00:03:24.19" />
                    <SPLIT distance="300" swimtime="00:04:06.33" />
                    <SPLIT distance="350" swimtime="00:04:47.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="James" lastname="Roberto Zoschke" birthdate="1976-02-08" gender="M" nation="BRA" license="312251" swrid="5688617" athleteid="9562" externalid="312251" level="DKMBANK">
              <RESULTS>
                <RESULT eventid="1123" points="399" swimtime="00:10:14.10" resultid="9563" heatid="10517" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                    <SPLIT distance="100" swimtime="00:01:12.86" />
                    <SPLIT distance="150" swimtime="00:01:51.49" />
                    <SPLIT distance="200" swimtime="00:02:30.18" />
                    <SPLIT distance="250" swimtime="00:03:09.07" />
                    <SPLIT distance="300" swimtime="00:03:48.31" />
                    <SPLIT distance="350" swimtime="00:04:27.38" />
                    <SPLIT distance="400" swimtime="00:05:06.68" />
                    <SPLIT distance="450" swimtime="00:05:45.33" />
                    <SPLIT distance="500" swimtime="00:06:24.58" />
                    <SPLIT distance="550" swimtime="00:07:03.24" />
                    <SPLIT distance="600" swimtime="00:07:42.23" />
                    <SPLIT distance="650" swimtime="00:08:20.91" />
                    <SPLIT distance="700" swimtime="00:08:59.80" />
                    <SPLIT distance="750" swimtime="00:09:37.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="424" swimtime="00:02:46.94" resultid="9564" heatid="10491" lane="0" entrytime="00:02:51.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.69" />
                    <SPLIT distance="100" swimtime="00:01:20.49" />
                    <SPLIT distance="150" swimtime="00:02:04.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="372" swimtime="00:20:10.20" resultid="9565" heatid="10637" lane="5" entrytime="00:19:49.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                    <SPLIT distance="100" swimtime="00:01:17.40" />
                    <SPLIT distance="150" swimtime="00:01:58.53" />
                    <SPLIT distance="200" swimtime="00:02:39.65" />
                    <SPLIT distance="250" swimtime="00:03:21.28" />
                    <SPLIT distance="300" swimtime="00:04:02.59" />
                    <SPLIT distance="350" swimtime="00:04:43.88" />
                    <SPLIT distance="400" swimtime="00:05:25.18" />
                    <SPLIT distance="450" swimtime="00:06:06.18" />
                    <SPLIT distance="500" swimtime="00:06:47.29" />
                    <SPLIT distance="550" swimtime="00:07:28.03" />
                    <SPLIT distance="600" swimtime="00:08:08.43" />
                    <SPLIT distance="650" swimtime="00:08:49.19" />
                    <SPLIT distance="700" swimtime="00:09:29.41" />
                    <SPLIT distance="750" swimtime="00:10:10.09" />
                    <SPLIT distance="800" swimtime="00:10:50.86" />
                    <SPLIT distance="850" swimtime="00:11:31.21" />
                    <SPLIT distance="900" swimtime="00:12:11.84" />
                    <SPLIT distance="950" swimtime="00:12:52.38" />
                    <SPLIT distance="1000" swimtime="00:13:32.88" />
                    <SPLIT distance="1050" swimtime="00:14:13.38" />
                    <SPLIT distance="1100" swimtime="00:14:53.74" />
                    <SPLIT distance="1150" swimtime="00:15:34.00" />
                    <SPLIT distance="1200" swimtime="00:16:14.31" />
                    <SPLIT distance="1250" swimtime="00:16:54.54" />
                    <SPLIT distance="1300" swimtime="00:17:34.70" />
                    <SPLIT distance="1350" swimtime="00:18:14.54" />
                    <SPLIT distance="1400" swimtime="00:18:53.82" />
                    <SPLIT distance="1450" swimtime="00:19:32.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="451" swimtime="00:01:14.15" resultid="9566" heatid="10598" lane="1" entrytime="00:01:13.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="403" swimtime="00:02:34.27" resultid="9567" heatid="10649" lane="4" entrytime="00:02:37.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                    <SPLIT distance="100" swimtime="00:01:13.74" />
                    <SPLIT distance="150" swimtime="00:01:58.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="429" swimtime="00:04:51.76" resultid="9568" heatid="10721" lane="2" entrytime="00:04:55.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                    <SPLIT distance="100" swimtime="00:01:09.94" />
                    <SPLIT distance="150" swimtime="00:01:47.15" />
                    <SPLIT distance="200" swimtime="00:02:24.28" />
                    <SPLIT distance="250" swimtime="00:03:01.65" />
                    <SPLIT distance="300" swimtime="00:03:38.92" />
                    <SPLIT distance="350" swimtime="00:04:16.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Victor Araujo" birthdate="2001-12-29" gender="M" nation="BRA" license="281163" swrid="5811241" athleteid="9511" externalid="281163" level="SMELJ | DK">
              <RESULTS>
                <RESULT eventid="1087" points="425" swimtime="00:02:46.86" resultid="9512" heatid="10487" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.32" />
                    <SPLIT distance="100" swimtime="00:01:21.34" />
                    <SPLIT distance="150" swimtime="00:02:05.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="706" swimtime="00:00:29.13" resultid="9513" heatid="10575" lane="4" entrytime="00:00:28.67" entrycourse="LCM" />
                <RESULT eventid="1235" points="585" swimtime="00:00:24.99" resultid="9514" heatid="10611" lane="5" />
                <RESULT eventid="1219" points="661" swimtime="00:01:05.28" resultid="9515" heatid="10599" lane="6" entrytime="00:01:04.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="501" swimtime="00:02:23.51" resultid="9516" heatid="10645" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.47" />
                    <SPLIT distance="100" swimtime="00:01:09.51" />
                    <SPLIT distance="150" swimtime="00:01:48.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="530" swimtime="00:01:03.74" resultid="9517" heatid="10733" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aline" lastname="Artigas" birthdate="1998-07-11" gender="F" nation="BRA" license="279942" athleteid="9500" externalid="279942">
              <RESULTS>
                <RESULT eventid="1095" points="276" swimtime="00:00:37.49" resultid="9501" heatid="10494" lane="5" />
                <RESULT eventid="1179" points="239" swimtime="00:00:46.93" resultid="9502" heatid="10561" lane="0" />
                <RESULT eventid="1147" points="319" swimtime="00:01:15.61" resultid="9503" heatid="10524" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="363" swimtime="00:00:33.07" resultid="9504" heatid="10600" lane="6" />
                <RESULT eventid="1297" points="272" swimtime="00:00:41.44" resultid="9505" heatid="10676" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Garcia Fraga" birthdate="2003-10-07" gender="M" nation="BRA" license="283467" swrid="5717265" athleteid="9536" externalid="283467" level="SMELJ | DK">
              <RESULTS>
                <RESULT eventid="1155" points="501" swimtime="00:00:58.41" resultid="9537" heatid="10550" lane="9" entrytime="00:00:57.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="420" swimtime="00:01:15.95" resultid="9538" heatid="10598" lane="9" entrytime="00:01:13.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" status="DNS" swimtime="00:00:00.00" resultid="9539" heatid="10682" lane="8" />
                <RESULT eventid="1273" points="495" swimtime="00:02:24.08" resultid="9540" heatid="10652" lane="9" entrytime="00:02:22.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.34" />
                    <SPLIT distance="100" swimtime="00:01:07.29" />
                    <SPLIT distance="150" swimtime="00:01:49.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="424" swimtime="00:01:05.82" resultid="9541" heatid="10709" lane="3" entrytime="00:01:04.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="461" swimtime="00:01:06.78" resultid="9542" heatid="10741" lane="9" entrytime="00:01:06.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Ocanha" birthdate="2005-06-21" gender="M" nation="BRA" license="313769" swrid="5600231" athleteid="9518" externalid="313769" level="SMELJ | DK">
              <RESULTS>
                <RESULT eventid="1103" points="496" swimtime="00:00:28.13" resultid="9519" heatid="10501" lane="1" />
                <RESULT eventid="1187" points="590" swimtime="00:00:30.93" resultid="9520" heatid="10575" lane="7" entrytime="00:00:30.60" entrycourse="LCM" />
                <RESULT eventid="1155" points="615" swimtime="00:00:54.54" resultid="9521" heatid="10551" lane="4" entrytime="00:00:54.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="605" swimtime="00:00:24.72" resultid="9522" heatid="10628" lane="1" entrytime="00:00:24.52" entrycourse="LCM" />
                <RESULT eventid="1305" points="459" swimtime="00:00:30.52" resultid="9523" heatid="10686" lane="4" entrytime="00:00:30.52" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isis" lastname="De Miranda" birthdate="2012-01-10" gender="F" nation="BRA" license="397278" swrid="5652886" athleteid="9603" externalid="397278" level="DKMBANK">
              <RESULTS>
                <RESULT eventid="1147" points="350" swimtime="00:01:13.34" resultid="9604" heatid="10527" lane="6" entrytime="00:01:15.42" entrycourse="LCM" />
                <RESULT eventid="1227" points="350" swimtime="00:00:33.50" resultid="9605" heatid="10602" lane="4" entrytime="00:00:34.96" entrycourse="LCM" />
                <RESULT eventid="1297" points="269" swimtime="00:00:41.60" resultid="9606" heatid="10677" lane="7" />
                <RESULT eventid="1281" points="322" swimtime="00:02:43.72" resultid="9607" heatid="10655" lane="8" entrytime="00:02:44.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                    <SPLIT distance="100" swimtime="00:01:18.24" />
                    <SPLIT distance="150" swimtime="00:02:01.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="277" swimtime="00:01:27.56" resultid="9608" heatid="10726" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Campesi" birthdate="2004-10-30" gender="M" nation="BRA" license="383112" swrid="5780365" athleteid="9581" externalid="383112" level="DKMBANK">
              <RESULTS>
                <RESULT eventid="1155" points="518" swimtime="00:00:57.76" resultid="9582" heatid="10549" lane="5" entrytime="00:00:57.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="576" swimtime="00:00:25.12" resultid="9583" heatid="10627" lane="8" entrytime="00:00:25.29" entrycourse="LCM" />
                <RESULT eventid="1289" points="357" swimtime="00:02:23.68" resultid="9584" heatid="10661" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                    <SPLIT distance="100" swimtime="00:01:04.87" />
                    <SPLIT distance="150" swimtime="00:01:42.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gilmar" lastname="Edson Schewtschik" birthdate="1982-07-17" gender="M" nation="BRA" license="053965" swrid="5810898" athleteid="9506" externalid="053965" level="DKMBANK">
              <RESULTS>
                <RESULT eventid="1187" points="340" swimtime="00:00:37.15" resultid="9507" heatid="10569" lane="1" />
                <RESULT eventid="1235" points="418" swimtime="00:00:27.95" resultid="9508" heatid="10622" lane="4" entrytime="00:00:27.90" entrycourse="LCM" />
                <RESULT eventid="1305" points="259" swimtime="00:00:36.93" resultid="9509" heatid="10682" lane="1" />
                <RESULT eventid="1289" points="335" swimtime="00:02:26.79" resultid="9510" heatid="10663" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                    <SPLIT distance="100" swimtime="00:01:06.36" />
                    <SPLIT distance="150" swimtime="00:01:45.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robson" lastname="Candido Dadalt" birthdate="1981-07-07" gender="M" nation="BRA" license="4637" swrid="5810812" athleteid="9591" externalid="4637" level="DKMBANK">
              <RESULTS>
                <RESULT eventid="1123" points="332" swimtime="00:10:52.63" resultid="9592" heatid="10517" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                    <SPLIT distance="100" swimtime="00:01:16.70" />
                    <SPLIT distance="150" swimtime="00:01:57.56" />
                    <SPLIT distance="200" swimtime="00:02:38.66" />
                    <SPLIT distance="250" swimtime="00:03:20.22" />
                    <SPLIT distance="300" swimtime="00:04:02.18" />
                    <SPLIT distance="350" swimtime="00:04:43.42" />
                    <SPLIT distance="400" swimtime="00:05:24.96" />
                    <SPLIT distance="450" swimtime="00:06:06.40" />
                    <SPLIT distance="500" swimtime="00:06:47.50" />
                    <SPLIT distance="550" swimtime="00:07:28.86" />
                    <SPLIT distance="600" swimtime="00:08:10.55" />
                    <SPLIT distance="650" swimtime="00:08:51.82" />
                    <SPLIT distance="700" swimtime="00:09:33.13" />
                    <SPLIT distance="750" swimtime="00:10:13.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="252" swimtime="00:02:56.96" resultid="9593" heatid="10475" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.86" />
                    <SPLIT distance="100" swimtime="00:01:26.12" />
                    <SPLIT distance="150" swimtime="00:02:11.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="341" swimtime="00:20:45.96" resultid="9594" heatid="10637" lane="8" entrytime="00:20:50.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                    <SPLIT distance="100" swimtime="00:01:16.06" />
                    <SPLIT distance="150" swimtime="00:01:56.77" />
                    <SPLIT distance="200" swimtime="00:02:37.73" />
                    <SPLIT distance="250" swimtime="00:03:19.05" />
                    <SPLIT distance="300" swimtime="00:04:00.23" />
                    <SPLIT distance="350" swimtime="00:04:41.83" />
                    <SPLIT distance="400" swimtime="00:05:23.30" />
                    <SPLIT distance="450" swimtime="00:06:05.13" />
                    <SPLIT distance="500" swimtime="00:06:46.28" />
                    <SPLIT distance="550" swimtime="00:07:27.79" />
                    <SPLIT distance="600" swimtime="00:08:09.24" />
                    <SPLIT distance="650" swimtime="00:08:50.54" />
                    <SPLIT distance="700" swimtime="00:09:32.77" />
                    <SPLIT distance="750" swimtime="00:10:14.63" />
                    <SPLIT distance="800" swimtime="00:10:56.65" />
                    <SPLIT distance="850" swimtime="00:11:38.86" />
                    <SPLIT distance="900" swimtime="00:12:21.46" />
                    <SPLIT distance="950" swimtime="00:13:04.12" />
                    <SPLIT distance="1000" swimtime="00:13:46.25" />
                    <SPLIT distance="1050" swimtime="00:14:28.64" />
                    <SPLIT distance="1100" swimtime="00:15:11.17" />
                    <SPLIT distance="1150" swimtime="00:15:53.29" />
                    <SPLIT distance="1200" swimtime="00:16:35.90" />
                    <SPLIT distance="1250" swimtime="00:17:18.43" />
                    <SPLIT distance="1300" swimtime="00:18:01.00" />
                    <SPLIT distance="1350" swimtime="00:18:43.55" />
                    <SPLIT distance="1400" swimtime="00:19:25.60" />
                    <SPLIT distance="1450" swimtime="00:20:07.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="306" swimtime="00:02:31.29" resultid="9595" heatid="10662" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                    <SPLIT distance="100" swimtime="00:01:11.63" />
                    <SPLIT distance="150" swimtime="00:01:51.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="348" swimtime="00:05:12.74" resultid="9596" heatid="10720" lane="1" entrytime="00:05:11.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                    <SPLIT distance="100" swimtime="00:01:14.90" />
                    <SPLIT distance="150" swimtime="00:01:54.39" />
                    <SPLIT distance="200" swimtime="00:02:34.19" />
                    <SPLIT distance="250" swimtime="00:03:13.78" />
                    <SPLIT distance="300" swimtime="00:03:53.79" />
                    <SPLIT distance="350" swimtime="00:04:33.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Angelo" lastname="De Queiroz" birthdate="2003-10-31" gender="M" nation="BRA" license="342814" swrid="5600149" athleteid="9549" externalid="342814" level="DKMBANK">
              <RESULTS>
                <RESULT eventid="1103" points="446" swimtime="00:00:29.14" resultid="9550" heatid="10507" lane="1" entrytime="00:00:28.60" entrycourse="LCM" />
                <RESULT eventid="1155" points="443" swimtime="00:01:00.86" resultid="9551" heatid="10547" lane="0" entrytime="00:01:02.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="395" swimtime="00:00:28.48" resultid="9552" heatid="10622" lane="0" entrytime="00:00:28.26" entrycourse="LCM" />
                <RESULT eventid="1305" points="374" swimtime="00:00:32.68" resultid="9553" heatid="10685" lane="3" entrytime="00:00:33.49" entrycourse="LCM" />
                <RESULT eventid="1341" points="402" swimtime="00:01:06.95" resultid="9554" heatid="10709" lane="7" entrytime="00:01:05.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="20" agetotalmax="-1" agetotalmin="-1" gender="M" name="WINNERS/DKMBANK &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1209" points="378" swimtime="00:09:38.79" resultid="9612" heatid="10582" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                    <SPLIT distance="100" swimtime="00:01:08.27" />
                    <SPLIT distance="150" swimtime="00:01:45.23" />
                    <SPLIT distance="200" swimtime="00:02:21.14" />
                    <SPLIT distance="250" swimtime="00:02:50.48" />
                    <SPLIT distance="300" swimtime="00:03:23.27" />
                    <SPLIT distance="350" swimtime="00:03:58.73" />
                    <SPLIT distance="400" swimtime="00:04:34.56" />
                    <SPLIT distance="450" swimtime="00:05:09.67" />
                    <SPLIT distance="500" swimtime="00:05:49.87" />
                    <SPLIT distance="550" swimtime="00:06:32.30" />
                    <SPLIT distance="600" swimtime="00:07:12.99" />
                    <SPLIT distance="650" swimtime="00:07:45.02" />
                    <SPLIT distance="700" swimtime="00:08:20.67" />
                    <SPLIT distance="750" swimtime="00:08:59.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9555" number="1" />
                    <RELAYPOSITION athleteid="9536" number="2" />
                    <RELAYPOSITION athleteid="9597" number="3" />
                    <RELAYPOSITION athleteid="9581" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="WINNERS/DKMBANK &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1331" points="527" swimtime="00:04:15.89" resultid="9613" heatid="10698" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                    <SPLIT distance="100" swimtime="00:01:05.38" />
                    <SPLIT distance="150" swimtime="00:01:37.25" />
                    <SPLIT distance="200" swimtime="00:02:16.45" />
                    <SPLIT distance="250" swimtime="00:02:46.49" />
                    <SPLIT distance="300" swimtime="00:03:19.98" />
                    <SPLIT distance="350" swimtime="00:03:46.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9536" number="1" />
                    <RELAYPOSITION athleteid="9518" number="2" />
                    <RELAYPOSITION athleteid="9569" number="3" />
                    <RELAYPOSITION athleteid="9543" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1399" points="574" swimtime="00:03:46.40" resultid="9614" heatid="10753" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.48" />
                    <SPLIT distance="100" swimtime="00:00:55.29" />
                    <SPLIT distance="150" swimtime="00:01:21.83" />
                    <SPLIT distance="200" swimtime="00:01:51.25" />
                    <SPLIT distance="250" swimtime="00:02:18.35" />
                    <SPLIT distance="300" swimtime="00:02:48.52" />
                    <SPLIT distance="350" swimtime="00:03:16.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9518" number="1" />
                    <RELAYPOSITION athleteid="9496" number="2" />
                    <RELAYPOSITION athleteid="9581" number="3" />
                    <RELAYPOSITION athleteid="9536" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="WINNERS/DKMBANK &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1331" points="425" swimtime="00:04:34.87" resultid="9616" heatid="10698" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                    <SPLIT distance="100" swimtime="00:01:09.44" />
                    <SPLIT distance="150" swimtime="00:01:45.82" />
                    <SPLIT distance="200" swimtime="00:02:25.62" />
                    <SPLIT distance="250" swimtime="00:02:57.99" />
                    <SPLIT distance="300" swimtime="00:03:34.96" />
                    <SPLIT distance="350" swimtime="00:04:04.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9496" number="1" />
                    <RELAYPOSITION athleteid="9562" number="2" />
                    <RELAYPOSITION athleteid="9549" number="3" />
                    <RELAYPOSITION athleteid="9581" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1399" points="499" swimtime="00:03:57.25" resultid="9617" heatid="10753" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.35" />
                    <SPLIT distance="100" swimtime="00:00:55.80" />
                    <SPLIT distance="150" swimtime="00:01:23.40" />
                    <SPLIT distance="200" swimtime="00:01:53.42" />
                    <SPLIT distance="250" swimtime="00:02:22.60" />
                    <SPLIT distance="300" swimtime="00:02:56.61" />
                    <SPLIT distance="350" swimtime="00:03:25.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9543" number="1" />
                    <RELAYPOSITION athleteid="9569" number="2" />
                    <RELAYPOSITION athleteid="9506" number="3" />
                    <RELAYPOSITION athleteid="9549" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="20" agetotalmax="-1" agetotalmin="-1" gender="F" name="WINNERS/DKMBANK &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1201" points="301" swimtime="00:11:22.55" resultid="9609" heatid="10578" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                    <SPLIT distance="100" swimtime="00:01:16.83" />
                    <SPLIT distance="150" swimtime="00:02:01.72" />
                    <SPLIT distance="200" swimtime="00:02:46.99" />
                    <SPLIT distance="250" swimtime="00:03:22.93" />
                    <SPLIT distance="300" swimtime="00:04:02.80" />
                    <SPLIT distance="350" swimtime="00:04:43.74" />
                    <SPLIT distance="450" swimtime="00:06:04.07" />
                    <SPLIT distance="500" swimtime="00:06:51.12" />
                    <SPLIT distance="550" swimtime="00:07:40.48" />
                    <SPLIT distance="650" swimtime="00:09:08.82" />
                    <SPLIT distance="700" swimtime="00:09:52.65" />
                    <SPLIT distance="750" swimtime="00:10:38.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9574" number="1" />
                    <RELAYPOSITION athleteid="9530" number="2" />
                    <RELAYPOSITION athleteid="9500" number="3" />
                    <RELAYPOSITION athleteid="9524" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="F" name="WINNERS/DKMBANK &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1321" points="289" swimtime="00:05:47.30" resultid="9610" heatid="10692" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.93" />
                    <SPLIT distance="100" swimtime="00:01:28.15" />
                    <SPLIT distance="150" swimtime="00:02:11.39" />
                    <SPLIT distance="200" swimtime="00:02:59.96" />
                    <SPLIT distance="250" swimtime="00:03:40.38" />
                    <SPLIT distance="350" swimtime="00:05:04.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9574" number="1" />
                    <RELAYPOSITION athleteid="9524" number="2" />
                    <RELAYPOSITION athleteid="9530" number="3" />
                    <RELAYPOSITION athleteid="9500" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1389" points="360" swimtime="00:04:52.21" resultid="9611" heatid="10747" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                    <SPLIT distance="100" swimtime="00:01:11.32" />
                    <SPLIT distance="150" swimtime="00:01:44.48" />
                    <SPLIT distance="200" swimtime="00:02:23.03" />
                    <SPLIT distance="250" swimtime="00:02:56.66" />
                    <SPLIT distance="300" swimtime="00:03:34.37" />
                    <SPLIT distance="350" swimtime="00:04:10.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9524" number="1" />
                    <RELAYPOSITION athleteid="9530" number="2" />
                    <RELAYPOSITION athleteid="9574" number="3" />
                    <RELAYPOSITION athleteid="9500" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="X" name="WINNERS/DKMBANK &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1247" points="416" swimtime="00:04:51.24" resultid="9615" heatid="10631" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                    <SPLIT distance="100" swimtime="00:01:07.35" />
                    <SPLIT distance="150" swimtime="00:01:49.91" />
                    <SPLIT distance="200" swimtime="00:02:37.14" />
                    <SPLIT distance="250" swimtime="00:03:06.58" />
                    <SPLIT distance="300" swimtime="00:03:39.73" />
                    <SPLIT distance="350" swimtime="00:04:12.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9536" number="1" />
                    <RELAYPOSITION athleteid="9530" number="2" />
                    <RELAYPOSITION athleteid="9569" number="3" />
                    <RELAYPOSITION athleteid="9524" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="X" name="WINNERS/DKMBANK &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1247" points="370" swimtime="00:05:02.62" resultid="9618" heatid="10631" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                    <SPLIT distance="100" swimtime="00:01:26.77" />
                    <SPLIT distance="150" swimtime="00:01:59.17" />
                    <SPLIT distance="200" swimtime="00:02:38.29" />
                    <SPLIT distance="250" swimtime="00:03:09.96" />
                    <SPLIT distance="300" swimtime="00:03:46.11" />
                    <SPLIT distance="350" swimtime="00:04:21.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9574" number="1" />
                    <RELAYPOSITION athleteid="9518" number="2" />
                    <RELAYPOSITION athleteid="9549" number="3" />
                    <RELAYPOSITION athleteid="9500" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="2864" nation="BRA" region="PR" clubid="6817" swrid="93756" name="Associacao De Pais E Amigos Da Natacao De Ponta Gr" shortname="Apan Ponta Grossa">
          <ATHLETES>
            <ATHLETE firstname="Augusto" lastname="Tramontin" birthdate="2011-11-29" gender="M" nation="BRA" license="399691" swrid="5652901" athleteid="6850" externalid="399691">
              <RESULTS>
                <RESULT eventid="1087" points="336" swimtime="00:03:00.42" resultid="6851" heatid="10489" lane="5" entrytime="00:03:02.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                    <SPLIT distance="100" swimtime="00:01:26.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="429" swimtime="00:00:34.39" resultid="6852" heatid="10573" lane="2" entrytime="00:00:35.99" entrycourse="LCM" />
                <RESULT eventid="1155" points="384" swimtime="00:01:03.79" resultid="6853" heatid="10546" lane="5" entrytime="00:01:02.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="411" swimtime="00:00:28.12" resultid="6854" heatid="10622" lane="6" entrytime="00:00:28.02" entrycourse="LCM" />
                <RESULT eventid="1219" points="377" swimtime="00:01:18.69" resultid="6855" heatid="10596" lane="0" entrytime="00:01:20.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="330" swimtime="00:00:34.06" resultid="6856" heatid="10685" lane="7" entrytime="00:00:35.37" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Pontes Mattioli" birthdate="2011-09-10" gender="F" nation="BRA" license="366914" swrid="5602572" athleteid="6870" externalid="366914">
              <RESULTS>
                <RESULT eventid="1095" points="355" swimtime="00:00:34.50" resultid="6871" heatid="10497" lane="8" entrytime="00:00:34.96" entrycourse="LCM" />
                <RESULT eventid="1063" points="333" swimtime="00:02:57.59" resultid="6872" heatid="10471" lane="0" entrytime="00:02:54.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.70" />
                    <SPLIT distance="100" swimtime="00:01:26.06" />
                    <SPLIT distance="150" swimtime="00:02:12.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="408" swimtime="00:01:09.71" resultid="6873" heatid="10530" lane="1" entrytime="00:01:08.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="429" swimtime="00:00:31.30" resultid="6874" heatid="10605" lane="9" entrytime="00:00:31.66" entrycourse="LCM" />
                <RESULT eventid="1297" points="355" swimtime="00:00:37.93" resultid="6875" heatid="10679" lane="2" entrytime="00:00:37.94" entrycourse="LCM" />
                <RESULT eventid="1365" points="349" swimtime="00:01:21.08" resultid="6876" heatid="10730" lane="1" entrytime="00:01:19.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Xavier Teixeira" birthdate="2011-09-22" gender="M" nation="BRA" license="415193" swrid="5762083" athleteid="6883" externalid="415193">
              <RESULTS>
                <RESULT eventid="1103" points="225" swimtime="00:00:36.61" resultid="6884" heatid="10501" lane="2" />
                <RESULT eventid="1187" points="139" swimtime="00:00:50.07" resultid="6885" heatid="10566" lane="4" />
                <RESULT eventid="1155" points="279" swimtime="00:01:10.94" resultid="6886" heatid="10541" lane="9" entrytime="00:01:12.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="272" swimtime="00:00:32.25" resultid="6887" heatid="10612" lane="1" />
                <RESULT eventid="1219" points="120" swimtime="00:01:55.09" resultid="6888" heatid="10591" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="174" swimtime="00:01:28.47" resultid="6889" heatid="10704" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Barbara" lastname="Campagnoli" birthdate="2009-04-13" gender="F" nation="BRA" license="366915" swrid="5600128" athleteid="6826" externalid="366915">
              <RESULTS>
                <RESULT eventid="1063" points="474" swimtime="00:02:37.83" resultid="6827" heatid="10473" lane="2" entrytime="00:02:35.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                    <SPLIT distance="100" swimtime="00:01:14.86" />
                    <SPLIT distance="150" swimtime="00:01:55.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="567" swimtime="00:01:02.44" resultid="6828" heatid="10534" lane="1" entrytime="00:01:03.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="590" swimtime="00:00:28.15" resultid="6829" heatid="10609" lane="7" entrytime="00:00:28.94" entrycourse="LCM" />
                <RESULT eventid="1297" points="539" swimtime="00:00:33.00" resultid="6830" heatid="10680" lane="6" entrytime="00:00:33.42" entrycourse="LCM" />
                <RESULT eventid="1365" points="456" swimtime="00:01:14.22" resultid="6831" heatid="10732" lane="6" entrytime="00:01:11.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Lievore" birthdate="2010-06-07" gender="F" nation="BRA" license="414856" swrid="5757092" athleteid="6861" externalid="414856">
              <RESULTS>
                <RESULT eventid="1147" points="339" swimtime="00:01:14.12" resultid="6862" heatid="10527" lane="4" entrytime="00:01:14.48" entrycourse="LCM" />
                <RESULT eventid="1227" points="331" swimtime="00:00:34.10" resultid="6863" heatid="10603" lane="8" entrytime="00:00:34.01" entrycourse="LCM" />
                <RESULT eventid="1297" points="265" swimtime="00:00:41.77" resultid="6864" heatid="10678" lane="3" entrytime="00:00:40.68" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Carraro Borges" birthdate="2009-05-11" gender="M" nation="BRA" license="345590" swrid="5622267" athleteid="6841" externalid="345590" level="SAGRADA FA">
              <RESULTS>
                <RESULT eventid="1123" points="426" swimtime="00:10:00.69" resultid="6842" heatid="10515" lane="4" entrytime="00:10:10.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                    <SPLIT distance="100" swimtime="00:01:06.23" />
                    <SPLIT distance="150" swimtime="00:01:43.12" />
                    <SPLIT distance="200" swimtime="00:02:21.21" />
                    <SPLIT distance="250" swimtime="00:02:59.27" />
                    <SPLIT distance="300" swimtime="00:03:38.02" />
                    <SPLIT distance="350" swimtime="00:04:17.36" />
                    <SPLIT distance="400" swimtime="00:04:56.85" />
                    <SPLIT distance="450" swimtime="00:05:35.93" />
                    <SPLIT distance="500" swimtime="00:06:14.88" />
                    <SPLIT distance="550" swimtime="00:06:54.16" />
                    <SPLIT distance="600" swimtime="00:07:32.73" />
                    <SPLIT distance="650" swimtime="00:08:10.76" />
                    <SPLIT distance="700" swimtime="00:08:49.19" />
                    <SPLIT distance="750" swimtime="00:09:26.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="423" swimtime="00:19:19.35" resultid="6843" heatid="10636" lane="1" entrytime="00:19:19.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                    <SPLIT distance="100" swimtime="00:01:10.31" />
                    <SPLIT distance="150" swimtime="00:01:48.35" />
                    <SPLIT distance="200" swimtime="00:02:27.49" />
                    <SPLIT distance="250" swimtime="00:03:05.76" />
                    <SPLIT distance="300" swimtime="00:03:45.09" />
                    <SPLIT distance="350" swimtime="00:04:24.88" />
                    <SPLIT distance="400" swimtime="00:05:04.75" />
                    <SPLIT distance="450" swimtime="00:05:44.94" />
                    <SPLIT distance="500" swimtime="00:06:24.16" />
                    <SPLIT distance="550" swimtime="00:07:04.90" />
                    <SPLIT distance="600" swimtime="00:07:46.01" />
                    <SPLIT distance="650" swimtime="00:08:26.15" />
                    <SPLIT distance="700" swimtime="00:09:05.30" />
                    <SPLIT distance="750" swimtime="00:09:44.36" />
                    <SPLIT distance="800" swimtime="00:10:23.79" />
                    <SPLIT distance="850" swimtime="00:11:02.43" />
                    <SPLIT distance="900" swimtime="00:11:41.49" />
                    <SPLIT distance="950" swimtime="00:12:20.14" />
                    <SPLIT distance="1000" swimtime="00:12:59.02" />
                    <SPLIT distance="1050" swimtime="00:13:37.35" />
                    <SPLIT distance="1100" swimtime="00:14:16.56" />
                    <SPLIT distance="1150" swimtime="00:14:55.19" />
                    <SPLIT distance="1200" swimtime="00:15:33.44" />
                    <SPLIT distance="1250" swimtime="00:16:11.24" />
                    <SPLIT distance="1300" swimtime="00:16:49.48" />
                    <SPLIT distance="1350" swimtime="00:17:27.25" />
                    <SPLIT distance="1400" swimtime="00:18:06.05" />
                    <SPLIT distance="1450" swimtime="00:18:43.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="417" swimtime="00:02:16.52" resultid="6844" heatid="10670" lane="6" entrytime="00:02:16.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.25" />
                    <SPLIT distance="100" swimtime="00:01:03.90" />
                    <SPLIT distance="150" swimtime="00:01:41.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="394" swimtime="00:05:00.10" resultid="6845" heatid="10722" lane="1" entrytime="00:04:47.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                    <SPLIT distance="100" swimtime="00:01:06.62" />
                    <SPLIT distance="150" swimtime="00:01:44.45" />
                    <SPLIT distance="200" swimtime="00:02:22.15" />
                    <SPLIT distance="250" swimtime="00:03:01.51" />
                    <SPLIT distance="300" swimtime="00:03:41.02" />
                    <SPLIT distance="350" swimtime="00:04:20.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Franca Berger" birthdate="2010-05-07" gender="F" nation="BRA" license="399692" swrid="5653290" athleteid="6865" externalid="399692">
              <RESULTS>
                <RESULT eventid="1095" points="205" swimtime="00:00:41.43" resultid="6866" heatid="10496" lane="0" entrytime="00:00:41.90" entrycourse="LCM" />
                <RESULT eventid="1147" points="287" swimtime="00:01:18.33" resultid="6867" heatid="10527" lane="0" entrytime="00:01:17.55" entrycourse="LCM" />
                <RESULT eventid="1227" points="309" swimtime="00:00:34.91" resultid="6868" heatid="10603" lane="0" entrytime="00:00:34.39" entrycourse="LCM" />
                <RESULT eventid="1211" points="248" swimtime="00:01:41.96" resultid="6869" heatid="10584" lane="1" entrytime="00:01:40.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yohan" lastname="Rigoni Moraes" birthdate="2002-04-03" gender="M" nation="BRA" license="272187" swrid="5600245" athleteid="6823" externalid="272187" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1187" points="691" swimtime="00:00:29.34" resultid="6824" heatid="10575" lane="5" entrytime="00:00:28.71" entrycourse="LCM" />
                <RESULT eventid="1219" points="624" swimtime="00:01:06.55" resultid="6825" heatid="10599" lane="1" entrytime="00:01:06.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Gueiber Montes" birthdate="2009-03-09" gender="M" nation="BRA" license="342154" swrid="5600179" athleteid="6818" externalid="342154">
              <RESULTS>
                <RESULT eventid="1155" points="625" swimtime="00:00:54.25" resultid="6819" heatid="10552" lane="8" entrytime="00:00:53.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="596" swimtime="00:00:24.84" resultid="6820" heatid="10628" lane="8" entrytime="00:00:24.54" entrycourse="LCM" />
                <RESULT eventid="1289" points="629" swimtime="00:01:58.99" resultid="6821" heatid="10674" lane="8" entrytime="00:01:59.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.05" />
                    <SPLIT distance="100" swimtime="00:00:56.73" />
                    <SPLIT distance="150" swimtime="00:01:27.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="593" swimtime="00:04:21.80" resultid="6822" heatid="10724" lane="8" entrytime="00:04:23.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                    <SPLIT distance="100" swimtime="00:01:01.40" />
                    <SPLIT distance="150" swimtime="00:01:35.13" />
                    <SPLIT distance="200" swimtime="00:02:08.55" />
                    <SPLIT distance="250" swimtime="00:02:42.86" />
                    <SPLIT distance="300" swimtime="00:03:16.90" />
                    <SPLIT distance="350" swimtime="00:03:49.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Brenda" lastname="Gabriele Carvalho" birthdate="2010-04-11" gender="F" nation="BRA" license="399557" swrid="5658060" athleteid="6857" externalid="399557">
              <RESULTS>
                <RESULT eventid="1079" points="278" swimtime="00:03:30.53" resultid="6858" heatid="10482" lane="2" entrytime="00:03:28.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.07" />
                    <SPLIT distance="100" swimtime="00:01:40.48" />
                    <SPLIT distance="150" swimtime="00:02:36.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="241" swimtime="00:00:46.85" resultid="6859" heatid="10562" lane="9" entrytime="00:00:48.36" entrycourse="LCM" />
                <RESULT eventid="1147" points="302" swimtime="00:01:17.04" resultid="6860" heatid="10527" lane="1" entrytime="00:01:16.26" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Sabedotti" birthdate="2011-04-20" gender="F" nation="BRA" license="390877" swrid="5602580" athleteid="6877" externalid="390877">
              <RESULTS>
                <RESULT eventid="1063" points="387" swimtime="00:02:48.86" resultid="6878" heatid="10471" lane="4" entrytime="00:02:50.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                    <SPLIT distance="100" swimtime="00:01:22.08" />
                    <SPLIT distance="150" swimtime="00:02:06.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="563" swimtime="00:01:02.62" resultid="6879" heatid="10533" lane="4" entrytime="00:01:04.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="512" swimtime="00:00:29.50" resultid="6880" heatid="10608" lane="9" entrytime="00:00:29.73" entrycourse="LCM" />
                <RESULT eventid="1281" points="532" swimtime="00:02:18.43" resultid="6881" heatid="10659" lane="2" entrytime="00:02:22.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                    <SPLIT distance="100" swimtime="00:01:06.18" />
                    <SPLIT distance="150" swimtime="00:01:42.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="405" swimtime="00:01:17.20" resultid="6882" heatid="10731" lane="9" entrytime="00:01:17.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Carolina Babiuki" birthdate="2007-02-06" gender="F" nation="BRA" license="316227" swrid="5600131" athleteid="6832" externalid="316227" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1227" points="528" swimtime="00:00:29.21" resultid="6833" heatid="10609" lane="6" entrytime="00:00:28.63" entrycourse="LCM" />
                <RESULT eventid="1297" points="520" swimtime="00:00:33.39" resultid="6834" heatid="10680" lane="3" entrytime="00:00:32.39" entrycourse="LCM" />
                <RESULT eventid="1365" points="453" swimtime="00:01:14.34" resultid="6835" heatid="10732" lane="2" entrytime="00:01:12.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yoseph" lastname="Rigoni Moraes" birthdate="2006-04-17" gender="M" nation="BRA" license="295182" swrid="5622302" athleteid="6846" externalid="295182" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1235" points="513" swimtime="00:00:26.12" resultid="6847" heatid="10625" lane="3" entrytime="00:00:26.11" entrycourse="LCM" />
                <RESULT eventid="1273" points="446" swimtime="00:02:29.16" resultid="6848" heatid="10650" lane="8" entrytime="00:02:33.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.50" />
                    <SPLIT distance="100" swimtime="00:01:09.52" />
                    <SPLIT distance="150" swimtime="00:01:53.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="386" swimtime="00:01:07.86" resultid="6849" heatid="10708" lane="3" entrytime="00:01:08.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Delinski" birthdate="2009-11-28" gender="F" nation="BRA" license="385190" swrid="5600150" athleteid="6836" externalid="385190">
              <RESULTS>
                <RESULT eventid="1079" points="327" swimtime="00:03:19.46" resultid="6837" heatid="10482" lane="4" entrytime="00:03:20.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.43" />
                    <SPLIT distance="100" swimtime="00:01:36.14" />
                    <SPLIT distance="150" swimtime="00:02:28.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="383" swimtime="00:00:40.14" resultid="6838" heatid="10564" lane="0" entrytime="00:00:40.10" entrycourse="LCM" />
                <RESULT eventid="1211" points="365" swimtime="00:01:29.68" resultid="6839" heatid="10587" lane="9" entrytime="00:01:26.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="356" swimtime="00:00:37.87" resultid="6840" heatid="10679" lane="5" entrytime="00:00:37.51" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="F" name="APAN/PONTA GROSSA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1387" points="408" swimtime="00:04:40.16" resultid="6890" heatid="10746" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                    <SPLIT distance="100" swimtime="00:01:01.78" />
                    <SPLIT distance="150" swimtime="00:01:35.80" />
                    <SPLIT distance="200" swimtime="00:02:13.06" />
                    <SPLIT distance="250" swimtime="00:02:47.21" />
                    <SPLIT distance="300" swimtime="00:03:28.36" />
                    <SPLIT distance="350" swimtime="00:04:02.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6826" number="1" />
                    <RELAYPOSITION athleteid="6836" number="2" />
                    <RELAYPOSITION athleteid="6865" number="3" />
                    <RELAYPOSITION athleteid="6861" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="APAN/PONTA GROSSA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1113" points="321" swimtime="00:05:17.50" resultid="6891" heatid="10510" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                    <SPLIT distance="100" swimtime="00:01:23.95" />
                    <SPLIT distance="150" swimtime="00:02:01.44" />
                    <SPLIT distance="200" swimtime="00:02:46.28" />
                    <SPLIT distance="250" swimtime="00:03:24.87" />
                    <SPLIT distance="300" swimtime="00:04:14.32" />
                    <SPLIT distance="350" swimtime="00:04:44.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6870" number="1" />
                    <RELAYPOSITION athleteid="6850" number="2" />
                    <RELAYPOSITION athleteid="6883" number="3" />
                    <RELAYPOSITION athleteid="6877" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="X" name="APAN/PONTA GROSSA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1245" points="436" swimtime="00:04:46.68" resultid="6892" heatid="10630" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="100" swimtime="00:01:14.32" />
                    <SPLIT distance="150" swimtime="00:01:54.72" />
                    <SPLIT distance="200" swimtime="00:02:42.36" />
                    <SPLIT distance="250" swimtime="00:03:11.95" />
                    <SPLIT distance="300" swimtime="00:03:46.80" />
                    <SPLIT distance="350" swimtime="00:04:14.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6826" number="1" />
                    <RELAYPOSITION athleteid="6836" number="2" />
                    <RELAYPOSITION athleteid="6818" number="3" />
                    <RELAYPOSITION athleteid="6841" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="2416" nation="BRA" region="PR" clubid="6893" swrid="93758" name="Apan/Maringá">
          <ATHLETES>
            <ATHLETE firstname="Gabriel" lastname="Antonio Mendes" birthdate="2008-12-04" gender="M" nation="BRA" license="366962" swrid="5196287" athleteid="6945" externalid="366962">
              <RESULTS>
                <RESULT eventid="1087" points="533" swimtime="00:02:34.71" resultid="6946" heatid="10492" lane="3" entrytime="00:02:31.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                    <SPLIT distance="100" swimtime="00:01:11.20" />
                    <SPLIT distance="150" swimtime="00:01:53.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="607" swimtime="00:00:30.64" resultid="6947" heatid="10575" lane="8" entrytime="00:00:30.92" entrycourse="LCM" />
                <RESULT eventid="1235" points="478" swimtime="00:00:26.73" resultid="6948" heatid="10611" lane="8" />
                <RESULT eventid="1219" points="563" swimtime="00:01:08.85" resultid="6949" heatid="10598" lane="4" entrytime="00:01:08.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="507" swimtime="00:00:29.52" resultid="6950" heatid="10686" lane="3" entrytime="00:00:30.89" entrycourse="LCM" />
                <RESULT eventid="1373" points="488" swimtime="00:01:05.51" resultid="6951" heatid="10741" lane="0" entrytime="00:01:06.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felype" lastname="Gongora Zago" birthdate="2011-09-14" gender="M" nation="BRA" license="392099" swrid="5603848" athleteid="6970" externalid="392099">
              <RESULTS>
                <RESULT eventid="1103" points="277" swimtime="00:00:34.13" resultid="6971" heatid="10503" lane="0" entrytime="00:00:37.06" entrycourse="LCM" />
                <RESULT eventid="1155" points="294" swimtime="00:01:09.76" resultid="6972" heatid="10539" lane="4" entrytime="00:01:14.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="297" swimtime="00:00:31.31" resultid="6973" heatid="10614" lane="4" entrytime="00:00:33.56" entrycourse="LCM" />
                <RESULT eventid="1341" points="159" swimtime="00:01:31.25" resultid="6974" heatid="10705" lane="9" entrytime="00:01:40.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Ayres" birthdate="2012-05-05" gender="M" nation="BRA" license="378035" swrid="5208079" athleteid="7033" externalid="378035">
              <RESULTS>
                <RESULT eventid="1071" points="341" swimtime="00:02:40.10" resultid="7034" heatid="10474" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                    <SPLIT distance="100" swimtime="00:01:17.27" />
                    <SPLIT distance="150" swimtime="00:02:00.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="300" swimtime="00:06:02.18" resultid="7035" heatid="10521" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.09" />
                    <SPLIT distance="100" swimtime="00:01:25.08" />
                    <SPLIT distance="150" swimtime="00:02:10.76" />
                    <SPLIT distance="200" swimtime="00:02:55.56" />
                    <SPLIT distance="250" swimtime="00:03:49.01" />
                    <SPLIT distance="300" swimtime="00:04:43.09" />
                    <SPLIT distance="350" swimtime="00:05:25.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="349" swimtime="00:00:33.44" resultid="7036" heatid="10685" lane="9" entrytime="00:00:35.83" entrycourse="LCM" />
                <RESULT eventid="1273" points="338" swimtime="00:02:43.64" resultid="7037" heatid="10645" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                    <SPLIT distance="100" swimtime="00:01:17.16" />
                    <SPLIT distance="150" swimtime="00:02:07.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="368" swimtime="00:05:06.99" resultid="7038" heatid="10720" lane="0" entrytime="00:05:15.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                    <SPLIT distance="100" swimtime="00:01:15.13" />
                    <SPLIT distance="150" swimtime="00:01:54.50" />
                    <SPLIT distance="200" swimtime="00:02:35.29" />
                    <SPLIT distance="250" swimtime="00:03:13.93" />
                    <SPLIT distance="300" swimtime="00:03:53.91" />
                    <SPLIT distance="350" swimtime="00:04:32.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Casavechia Carraro" birthdate="2009-07-28" gender="M" nation="BRA" license="368150" swrid="5384752" athleteid="6894" externalid="368150">
              <RESULTS>
                <RESULT eventid="1103" points="656" swimtime="00:00:25.62" resultid="6895" heatid="10508" lane="2" entrytime="00:00:26.75" entrycourse="LCM" />
                <RESULT eventid="1155" points="688" swimtime="00:00:52.55" resultid="6896" heatid="10552" lane="3" entrytime="00:00:52.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="606" swimtime="00:00:24.70" resultid="6897" heatid="10627" lane="4" entrytime="00:00:24.82" entrycourse="LCM" />
                <RESULT eventid="1289" points="648" swimtime="00:01:57.84" resultid="6898" heatid="10674" lane="6" entrytime="00:01:57.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.30" />
                    <SPLIT distance="100" swimtime="00:00:57.88" />
                    <SPLIT distance="150" swimtime="00:01:27.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="647" swimtime="00:00:57.15" resultid="6899" heatid="10711" lane="4" entrytime="00:00:57.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Garcia Cavalcante" birthdate="2011-11-21" gender="M" nation="BRA" license="378200" swrid="5603840" athleteid="6925" externalid="378200">
              <RESULTS>
                <RESULT eventid="1087" points="350" swimtime="00:02:58.02" resultid="6926" heatid="10489" lane="1" entrytime="00:03:10.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                    <SPLIT distance="100" swimtime="00:01:27.58" />
                    <SPLIT distance="150" swimtime="00:02:15.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="342" swimtime="00:00:37.08" resultid="6927" heatid="10572" lane="2" entrytime="00:00:39.38" entrycourse="LCM" />
                <RESULT eventid="1219" points="363" swimtime="00:01:19.68" resultid="6928" heatid="10594" lane="6" entrytime="00:01:26.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="308" swimtime="00:02:48.72" resultid="6929" heatid="10647" lane="0" entrytime="00:03:05.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.77" />
                    <SPLIT distance="100" swimtime="00:01:23.22" />
                    <SPLIT distance="150" swimtime="00:02:11.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Marques Picolo Vinha" birthdate="2010-07-01" gender="M" nation="BRA" license="366990" swrid="5603869" athleteid="6964" externalid="366990">
              <RESULTS>
                <RESULT eventid="1155" points="414" swimtime="00:01:02.25" resultid="6965" heatid="10545" lane="0" entrytime="00:01:05.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="386" swimtime="00:00:28.70" resultid="6966" heatid="10620" lane="2" entrytime="00:00:29.43" entrycourse="LCM" />
                <RESULT eventid="1305" points="327" swimtime="00:00:34.16" resultid="6967" heatid="10682" lane="3" />
                <RESULT eventid="1289" points="357" swimtime="00:02:23.67" resultid="6968" heatid="10667" lane="5" entrytime="00:02:27.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:08.19" />
                    <SPLIT distance="150" swimtime="00:01:47.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="308" swimtime="00:01:16.39" resultid="6969" heatid="10737" lane="8" entrytime="00:01:18.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Diogo" lastname="Sanchez" birthdate="2012-11-29" gender="M" nation="BRA" license="370658" swrid="5603906" athleteid="6930" externalid="370658">
              <RESULTS>
                <RESULT eventid="1087" points="233" swimtime="00:03:23.78" resultid="6931" heatid="10487" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.00" />
                    <SPLIT distance="100" swimtime="00:01:39.96" />
                    <SPLIT distance="150" swimtime="00:02:34.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="235" swimtime="00:00:42.01" resultid="6932" heatid="10569" lane="8" />
                <RESULT eventid="1219" points="219" swimtime="00:01:34.23" resultid="6933" heatid="10591" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Chaim" birthdate="2011-05-29" gender="F" nation="BRA" license="370662" swrid="5409721" athleteid="7004" externalid="370662">
              <RESULTS>
                <RESULT eventid="1063" points="273" swimtime="00:03:09.69" resultid="7005" heatid="10469" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="364" swimtime="00:01:12.42" resultid="7006" heatid="10527" lane="5" entrytime="00:01:14.73" entrycourse="LCM" />
                <RESULT eventid="1227" points="369" swimtime="00:00:32.89" resultid="7007" heatid="10603" lane="2" entrytime="00:00:33.11" entrycourse="LCM" />
                <RESULT eventid="1281" points="317" swimtime="00:02:44.48" resultid="7008" heatid="10654" lane="5" entrytime="00:02:48.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.36" />
                    <SPLIT distance="100" swimtime="00:01:18.53" />
                    <SPLIT distance="150" swimtime="00:02:02.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="262" swimtime="00:01:29.18" resultid="7009" heatid="10727" lane="3" entrytime="00:01:31.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Mochiutti Carneiro" birthdate="2010-04-22" gender="F" nation="BRA" license="370670" swrid="5588817" athleteid="6998" externalid="370670">
              <RESULTS>
                <RESULT eventid="1095" points="392" swimtime="00:00:33.38" resultid="6999" heatid="10498" lane="0" entrytime="00:00:33.06" entrycourse="LCM" />
                <RESULT eventid="1147" points="486" swimtime="00:01:05.73" resultid="7000" heatid="10533" lane="6" entrytime="00:01:04.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="435" swimtime="00:00:31.16" resultid="7001" heatid="10607" lane="5" entrytime="00:00:29.92" entrycourse="LCM" />
                <RESULT eventid="1281" points="477" swimtime="00:02:23.63" resultid="7002" heatid="10658" lane="4" entrytime="00:02:24.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                    <SPLIT distance="100" swimtime="00:01:09.97" />
                    <SPLIT distance="150" swimtime="00:01:47.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="365" swimtime="00:01:17.17" resultid="7003" heatid="10702" lane="0" entrytime="00:01:13.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Passafaro" birthdate="2009-02-01" gender="F" nation="BRA" license="370673" swrid="5603885" athleteid="6940" externalid="370673">
              <RESULTS>
                <RESULT eventid="1095" points="388" swimtime="00:00:33.47" resultid="6941" heatid="10497" lane="6" entrytime="00:00:34.38" entrycourse="LCM" />
                <RESULT eventid="1147" points="386" swimtime="00:01:10.96" resultid="6942" heatid="10528" lane="9" entrytime="00:01:14.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="421" swimtime="00:00:31.49" resultid="6943" heatid="10606" lane="0" entrytime="00:00:31.15" entrycourse="LCM" />
                <RESULT eventid="1333" points="333" swimtime="00:01:19.59" resultid="6944" heatid="10700" lane="6" entrytime="00:01:29.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Pacheco" birthdate="2006-12-20" gender="M" nation="BRA" license="336850" swrid="5603854" athleteid="6934" externalid="336850">
              <RESULTS>
                <RESULT eventid="1103" points="479" swimtime="00:00:28.45" resultid="6935" heatid="10507" lane="3" entrytime="00:00:28.20" entrycourse="LCM" />
                <RESULT eventid="1171" points="399" swimtime="00:02:29.81" resultid="6936" heatid="10555" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.15" />
                    <SPLIT distance="100" swimtime="00:01:06.05" />
                    <SPLIT distance="150" swimtime="00:01:46.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="481" swimtime="00:00:26.68" resultid="6937" heatid="10625" lane="1" entrytime="00:00:26.78" entrycourse="LCM" />
                <RESULT eventid="1273" points="476" swimtime="00:02:25.94" resultid="6938" heatid="10650" lane="7" entrytime="00:02:33.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                    <SPLIT distance="100" swimtime="00:01:07.09" />
                    <SPLIT distance="150" swimtime="00:01:53.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="481" swimtime="00:01:03.07" resultid="6939" heatid="10710" lane="8" entrytime="00:01:03.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Corsine Ferreira" birthdate="2010-03-10" gender="F" nation="BRA" license="353591" swrid="5588608" athleteid="6993" externalid="353591">
              <RESULTS>
                <RESULT eventid="1063" points="315" swimtime="00:03:00.97" resultid="6994" heatid="10472" lane="9" entrytime="00:02:49.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                    <SPLIT distance="100" swimtime="00:01:25.39" />
                    <SPLIT distance="150" swimtime="00:02:13.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="277" swimtime="00:00:44.69" resultid="6995" heatid="10564" lane="9" entrytime="00:00:40.21" entrycourse="LCM" />
                <RESULT eventid="1297" points="371" swimtime="00:00:37.38" resultid="6996" heatid="10680" lane="1" entrytime="00:00:35.40" entrycourse="LCM" />
                <RESULT eventid="1365" points="325" swimtime="00:01:23.03" resultid="6997" heatid="10730" lane="4" entrytime="00:01:17.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edgar" lastname="Romero" birthdate="2011-05-12" gender="M" nation="BRA" license="413920" athleteid="7061" externalid="413920">
              <RESULTS>
                <RESULT eventid="1155" points="353" swimtime="00:01:05.64" resultid="7062" heatid="10535" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="363" swimtime="00:00:29.29" resultid="7063" heatid="10613" lane="8" />
                <RESULT eventid="1289" points="312" swimtime="00:02:30.30" resultid="7064" heatid="10661" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                    <SPLIT distance="100" swimtime="00:01:10.18" />
                    <SPLIT distance="150" swimtime="00:01:51.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="281" swimtime="00:05:35.61" resultid="7065" heatid="10717" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                    <SPLIT distance="100" swimtime="00:01:13.60" />
                    <SPLIT distance="150" swimtime="00:01:57.11" />
                    <SPLIT distance="200" swimtime="00:02:41.16" />
                    <SPLIT distance="250" swimtime="00:03:25.95" />
                    <SPLIT distance="300" swimtime="00:04:10.35" />
                    <SPLIT distance="350" swimtime="00:04:55.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hammon" lastname="Henrique Costa" birthdate="2008-09-19" gender="M" nation="BRA" license="408703" swrid="5726000" athleteid="7056" externalid="408703">
              <RESULTS>
                <RESULT eventid="1187" points="416" swimtime="00:00:34.76" resultid="7057" heatid="10567" lane="7" />
                <RESULT eventid="1155" points="381" swimtime="00:01:03.95" resultid="7058" heatid="10537" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="401" swimtime="00:00:28.35" resultid="7059" heatid="10611" lane="6" />
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 9:24)" eventid="1219" status="DSQ" swimtime="00:01:20.47" resultid="7060" heatid="10590" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lara" lastname="Constantino" birthdate="2012-06-02" gender="F" nation="BRA" license="382208" swrid="5420069" athleteid="7045" externalid="382208">
              <RESULTS>
                <RESULT eventid="1079" points="335" swimtime="00:03:17.89" resultid="7046" heatid="10481" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.89" />
                    <SPLIT distance="100" swimtime="00:01:38.39" />
                    <SPLIT distance="150" swimtime="00:02:28.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="337" swimtime="00:00:41.90" resultid="7047" heatid="10563" lane="9" entrytime="00:00:42.89" entrycourse="LCM" />
                <RESULT eventid="1211" points="325" swimtime="00:01:33.26" resultid="7048" heatid="10584" lane="3" entrytime="00:01:37.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="270" swimtime="00:03:14.92" resultid="7049" heatid="10639" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.84" />
                    <SPLIT distance="100" swimtime="00:01:41.07" />
                    <SPLIT distance="150" swimtime="00:02:32.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Batista Sanchez" birthdate="2009-05-22" gender="M" nation="BRA" license="370668" swrid="5255779" athleteid="6913" externalid="370668">
              <RESULTS>
                <RESULT eventid="1087" points="418" swimtime="00:02:47.77" resultid="6914" heatid="10491" lane="5" entrytime="00:02:45.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                    <SPLIT distance="100" swimtime="00:01:18.28" />
                    <SPLIT distance="150" swimtime="00:02:03.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="427" swimtime="00:00:34.45" resultid="6915" heatid="10574" lane="6" entrytime="00:00:33.80" entrycourse="LCM" />
                <RESULT eventid="1235" points="381" swimtime="00:00:28.82" resultid="6916" heatid="10612" lane="8" />
                <RESULT eventid="1219" points="436" swimtime="00:01:14.98" resultid="6917" heatid="10597" lane="3" entrytime="00:01:14.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="346" swimtime="00:01:10.41" resultid="6918" heatid="10708" lane="0" entrytime="00:01:10.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Pavão" birthdate="2012-04-04" gender="F" nation="BRA" license="377259" swrid="5603888" athleteid="7022" externalid="377259">
              <RESULTS>
                <RESULT eventid="1063" points="320" swimtime="00:02:59.85" resultid="7023" heatid="10469" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="342" swimtime="00:01:13.89" resultid="7024" heatid="10526" lane="5" entrytime="00:01:19.28" entrycourse="LCM" />
                <RESULT eventid="1297" points="349" swimtime="00:00:38.15" resultid="7025" heatid="10678" lane="5" entrytime="00:00:40.09" entrycourse="LCM" />
                <RESULT eventid="1365" points="321" swimtime="00:01:23.36" resultid="7026" heatid="10728" lane="3" entrytime="00:01:27.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathan" lastname="Novak Pinho" birthdate="2012-11-14" gender="M" nation="BRA" license="378199" swrid="5603879" athleteid="7039" externalid="378199">
              <RESULTS>
                <RESULT eventid="1071" points="225" swimtime="00:03:03.83" resultid="7040" heatid="10474" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.50" />
                    <SPLIT distance="100" swimtime="00:01:29.15" />
                    <SPLIT distance="150" swimtime="00:02:17.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="270" swimtime="00:01:11.74" resultid="7041" heatid="10539" lane="3" entrytime="00:01:14.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="268" swimtime="00:00:32.42" resultid="7042" heatid="10614" lane="8" entrytime="00:00:35.36" entrycourse="LCM" />
                <RESULT eventid="1289" points="255" swimtime="00:02:40.72" resultid="7043" heatid="10665" lane="3" entrytime="00:02:44.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.95" />
                    <SPLIT distance="100" swimtime="00:01:15.72" />
                    <SPLIT distance="150" swimtime="00:01:57.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="256" swimtime="00:05:46.25" resultid="7044" heatid="10719" lane="0" entrytime="00:05:54.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                    <SPLIT distance="100" swimtime="00:01:18.59" />
                    <SPLIT distance="150" swimtime="00:02:01.76" />
                    <SPLIT distance="200" swimtime="00:02:46.69" />
                    <SPLIT distance="250" swimtime="00:03:31.11" />
                    <SPLIT distance="300" swimtime="00:04:17.38" />
                    <SPLIT distance="350" swimtime="00:05:01.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietro" lastname="Nabas De Assis" birthdate="2011-07-09" gender="M" nation="BRA" license="366968" swrid="5603878" athleteid="6981" externalid="366968">
              <RESULTS>
                <RESULT eventid="1087" points="309" swimtime="00:03:05.46" resultid="6982" heatid="10490" lane="2" entrytime="00:02:56.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.74" />
                    <SPLIT distance="100" swimtime="00:01:28.85" />
                    <SPLIT distance="150" swimtime="00:02:17.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="421" swimtime="00:00:34.62" resultid="6983" heatid="10573" lane="5" entrytime="00:00:35.74" entrycourse="LCM" />
                <RESULT eventid="1219" points="376" swimtime="00:01:18.79" resultid="6984" heatid="10597" lane="8" entrytime="00:01:18.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="316" swimtime="00:02:29.71" resultid="6985" heatid="10667" lane="9" entrytime="00:02:31.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                    <SPLIT distance="100" swimtime="00:01:10.72" />
                    <SPLIT distance="150" swimtime="00:01:50.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="340" swimtime="00:05:15.25" resultid="6986" heatid="10717" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                    <SPLIT distance="100" swimtime="00:01:13.42" />
                    <SPLIT distance="150" swimtime="00:01:53.89" />
                    <SPLIT distance="200" swimtime="00:02:35.15" />
                    <SPLIT distance="250" swimtime="00:03:16.15" />
                    <SPLIT distance="300" swimtime="00:03:57.23" />
                    <SPLIT distance="350" swimtime="00:04:37.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniela" lastname="Inoue" birthdate="2008-10-31" gender="F" nation="BRA" license="378348" swrid="5603856" athleteid="6958" externalid="378348">
              <RESULTS>
                <RESULT eventid="1063" points="254" swimtime="00:03:14.30" resultid="6959" heatid="10469" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="376" swimtime="00:01:11.64" resultid="6960" heatid="10529" lane="7" entrytime="00:01:10.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="372" swimtime="00:00:32.80" resultid="6961" heatid="10605" lane="4" entrytime="00:00:31.26" entrycourse="LCM" />
                <RESULT eventid="1297" points="308" swimtime="00:00:39.74" resultid="6962" heatid="10679" lane="7" entrytime="00:00:37.95" entrycourse="LCM" />
                <RESULT eventid="1365" points="280" swimtime="00:01:27.26" resultid="6963" heatid="10729" lane="8" entrytime="00:01:24.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Otavio Costa" birthdate="2009-01-28" gender="M" nation="BRA" license="370666" swrid="5603881" athleteid="6975" externalid="370666">
              <RESULTS>
                <RESULT eventid="1087" points="296" swimtime="00:03:08.26" resultid="6976" heatid="10489" lane="0" entrytime="00:03:12.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.81" />
                    <SPLIT distance="100" swimtime="00:01:29.28" />
                    <SPLIT distance="150" swimtime="00:02:18.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="266" swimtime="00:00:40.32" resultid="6977" heatid="10572" lane="1" entrytime="00:00:39.54" entrycourse="LCM" />
                <RESULT eventid="1155" points="340" swimtime="00:01:06.47" resultid="6978" heatid="10535" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="266" swimtime="00:01:28.34" resultid="6979" heatid="10594" lane="8" entrytime="00:01:27.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="326" swimtime="00:05:19.68" resultid="6980" heatid="10718" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                    <SPLIT distance="100" swimtime="00:01:15.54" />
                    <SPLIT distance="150" swimtime="00:01:56.16" />
                    <SPLIT distance="200" swimtime="00:02:37.83" />
                    <SPLIT distance="250" swimtime="00:03:19.41" />
                    <SPLIT distance="300" swimtime="00:04:00.99" />
                    <SPLIT distance="350" swimtime="00:04:42.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raphael" lastname="Piai Pellegrini" birthdate="2012-03-24" gender="M" nation="BRA" license="377261" swrid="5603894" athleteid="7027" externalid="377261">
              <RESULTS>
                <RESULT eventid="1103" points="394" swimtime="00:00:30.37" resultid="7028" heatid="10504" lane="2" entrytime="00:00:33.69" entrycourse="LCM" />
                <RESULT eventid="1155" points="443" swimtime="00:01:00.86" resultid="7029" heatid="10543" lane="3" entrytime="00:01:06.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="445" swimtime="00:00:27.37" resultid="7030" heatid="10793" lane="5" entrytime="00:00:29.40" entrycourse="LCM" />
                <RESULT eventid="1289" points="363" swimtime="00:02:22.91" resultid="7031" heatid="10663" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.47" />
                    <SPLIT distance="100" swimtime="00:01:08.89" />
                    <SPLIT distance="150" swimtime="00:01:48.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="316" swimtime="00:01:12.57" resultid="7032" heatid="10706" lane="0" entrytime="00:01:19.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wellington" lastname="De Lima" birthdate="2008-03-01" gender="M" nation="BRA" license="370024" swrid="5470912" athleteid="6906" externalid="370024">
              <RESULTS>
                <RESULT eventid="1103" points="460" swimtime="00:00:28.84" resultid="6907" heatid="10507" lane="0" entrytime="00:00:28.83" entrycourse="LCM" />
                <RESULT eventid="1155" points="553" swimtime="00:00:56.51" resultid="6908" heatid="10550" lane="1" entrytime="00:00:57.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="500" swimtime="00:00:26.33" resultid="6909" heatid="10625" lane="5" entrytime="00:00:26.09" entrycourse="LCM" />
                <RESULT eventid="1305" points="467" swimtime="00:00:30.34" resultid="6910" heatid="10686" lane="6" entrytime="00:00:31.23" entrycourse="LCM" />
                <RESULT eventid="1289" points="518" swimtime="00:02:07.00" resultid="6911" heatid="10671" lane="2" entrytime="00:02:13.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.31" />
                    <SPLIT distance="100" swimtime="00:01:00.06" />
                    <SPLIT distance="150" swimtime="00:01:33.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="430" swimtime="00:01:08.36" resultid="6912" heatid="10739" lane="6" entrytime="00:01:10.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Pacheco" birthdate="2012-10-03" gender="M" nation="BRA" license="370663" swrid="5603883" athleteid="7016" externalid="370663">
              <RESULTS>
                <RESULT eventid="1103" points="292" swimtime="00:00:33.54" resultid="7017" heatid="10504" lane="9" entrytime="00:00:34.74" entrycourse="LCM" />
                <RESULT eventid="1187" points="279" swimtime="00:00:39.68" resultid="7018" heatid="10568" lane="6" />
                <RESULT eventid="1155" points="288" swimtime="00:01:10.20" resultid="7019" heatid="10541" lane="1" entrytime="00:01:11.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="313" swimtime="00:00:30.78" resultid="7020" heatid="10793" lane="3" entrytime="00:00:31.70" entrycourse="LCM" />
                <RESULT eventid="1341" points="190" swimtime="00:01:26.01" resultid="7021" heatid="10703" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Ghelere" birthdate="2011-04-03" gender="F" nation="BRA" license="368146" swrid="5603843" athleteid="7010" externalid="368146">
              <RESULTS>
                <RESULT eventid="1095" points="349" swimtime="00:00:34.68" resultid="7011" heatid="10496" lane="3" entrytime="00:00:36.66" entrycourse="LCM" />
                <RESULT eventid="1147" points="338" swimtime="00:01:14.19" resultid="7012" heatid="10528" lane="7" entrytime="00:01:13.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="348" swimtime="00:00:33.55" resultid="7013" heatid="10603" lane="1" entrytime="00:00:33.91" entrycourse="LCM" />
                <RESULT eventid="1297" points="335" swimtime="00:00:38.67" resultid="7014" heatid="10677" lane="1" />
                <RESULT eventid="1365" points="308" swimtime="00:01:24.59" resultid="7015" heatid="10728" lane="4" entrytime="00:01:26.22" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Quental De Meireles" birthdate="2008-11-20" gender="M" nation="BRA" license="392103" swrid="5603898" athleteid="6987" externalid="392103">
              <RESULTS>
                <RESULT eventid="1103" points="425" swimtime="00:00:29.62" resultid="6988" heatid="10506" lane="5" entrytime="00:00:29.96" entrycourse="LCM" />
                <RESULT eventid="1187" points="386" swimtime="00:00:35.63" resultid="6989" heatid="10573" lane="6" entrytime="00:00:35.96" entrycourse="LCM" />
                <RESULT eventid="1235" points="372" swimtime="00:00:29.06" resultid="6990" heatid="10621" lane="7" entrytime="00:00:28.67" entrycourse="LCM" />
                <RESULT eventid="1289" points="393" swimtime="00:02:19.16" resultid="6991" heatid="10662" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.36" />
                    <SPLIT distance="100" swimtime="00:01:04.44" />
                    <SPLIT distance="150" swimtime="00:01:41.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="421" swimtime="00:01:05.96" resultid="6992" heatid="10708" lane="6" entrytime="00:01:08.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Muniz" birthdate="2012-09-03" gender="M" nation="BRA" license="392106" swrid="5603877" athleteid="7050" externalid="392106">
              <RESULTS>
                <RESULT eventid="1071" points="178" swimtime="00:03:18.69" resultid="7051" heatid="10474" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.90" />
                    <SPLIT distance="100" swimtime="00:01:36.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="263" swimtime="00:01:12.38" resultid="7052" heatid="10538" lane="1" entrytime="00:01:23.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="254" swimtime="00:00:33.01" resultid="7053" heatid="10613" lane="5" entrytime="00:00:36.26" entrycourse="LCM" />
                <RESULT eventid="1305" points="174" swimtime="00:00:42.16" resultid="7054" heatid="10683" lane="3" entrytime="00:00:48.29" entrycourse="LCM" />
                <RESULT eventid="1373" points="180" swimtime="00:01:31.37" resultid="7055" heatid="10735" lane="6" entrytime="00:01:54.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Biason Santana" birthdate="2009-01-21" gender="M" nation="BRA" license="366969" swrid="5317765" athleteid="6952" externalid="366969">
              <RESULTS>
                <RESULT eventid="1103" points="486" swimtime="00:00:28.32" resultid="6953" heatid="10507" lane="5" entrytime="00:00:27.76" entrycourse="LCM" />
                <RESULT eventid="1171" points="414" swimtime="00:02:27.99" resultid="6954" heatid="10557" lane="5" entrytime="00:02:28.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                    <SPLIT distance="100" swimtime="00:01:09.13" />
                    <SPLIT distance="150" swimtime="00:01:48.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="441" swimtime="00:00:27.46" resultid="6955" heatid="10624" lane="3" entrytime="00:00:27.04" entrycourse="LCM" />
                <RESULT eventid="1305" points="338" swimtime="00:00:33.79" resultid="6956" heatid="10682" lane="9" />
                <RESULT eventid="1341" points="493" swimtime="00:01:02.58" resultid="6957" heatid="10710" lane="7" entrytime="00:01:02.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Garcia Cavalcante" birthdate="2008-08-11" gender="M" nation="BRA" license="369676" swrid="5603841" athleteid="6919" externalid="369676">
              <RESULTS>
                <RESULT eventid="1087" points="374" swimtime="00:02:54.12" resultid="6920" heatid="10491" lane="6" entrytime="00:02:47.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.02" />
                    <SPLIT distance="100" swimtime="00:01:22.48" />
                    <SPLIT distance="150" swimtime="00:02:08.02" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 19:36)" eventid="1187" status="DSQ" swimtime="00:00:37.05" resultid="6921" heatid="10574" lane="0" entrytime="00:00:35.06" entrycourse="LCM" />
                <RESULT eventid="1219" status="DNS" swimtime="00:00:00.00" resultid="6922" heatid="10597" lane="7" entrytime="00:01:17.42" entrycourse="LCM" />
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 16:47)" eventid="1273" status="DSQ" swimtime="00:02:36.32" resultid="6923" heatid="10649" lane="5" entrytime="00:02:37.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                    <SPLIT distance="100" swimtime="00:01:14.53" />
                    <SPLIT distance="150" swimtime="00:01:59.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="393" swimtime="00:05:00.34" resultid="6924" heatid="10721" lane="0" entrytime="00:04:58.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                    <SPLIT distance="100" swimtime="00:01:10.45" />
                    <SPLIT distance="150" swimtime="00:01:48.75" />
                    <SPLIT distance="200" swimtime="00:02:27.37" />
                    <SPLIT distance="250" swimtime="00:03:04.70" />
                    <SPLIT distance="300" swimtime="00:03:43.43" />
                    <SPLIT distance="350" swimtime="00:04:21.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Campelo" birthdate="2011-09-12" gender="M" nation="BRA" license="366963" swrid="5588742" athleteid="6900" externalid="366963">
              <RESULTS>
                <RESULT eventid="1103" points="455" swimtime="00:00:28.94" resultid="6901" heatid="10506" lane="3" entrytime="00:00:30.16" entrycourse="LCM" />
                <RESULT eventid="1155" points="487" swimtime="00:00:58.97" resultid="6902" heatid="10550" lane="0" entrytime="00:00:57.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="526" swimtime="00:00:25.90" resultid="6903" heatid="10627" lane="9" entrytime="00:00:25.52" entrycourse="LCM" />
                <RESULT eventid="1289" points="442" swimtime="00:02:13.88" resultid="6904" heatid="10670" lane="5" entrytime="00:02:16.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.05" />
                    <SPLIT distance="100" swimtime="00:01:02.62" />
                    <SPLIT distance="150" swimtime="00:01:38.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="383" swimtime="00:01:08.06" resultid="6905" heatid="10708" lane="9" entrytime="00:01:10.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1331" points="493" swimtime="00:04:21.72" resultid="7068" heatid="10698" lane="5" entrytime="00:04:13.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                    <SPLIT distance="100" swimtime="00:01:10.88" />
                    <SPLIT distance="150" swimtime="00:01:41.89" />
                    <SPLIT distance="200" swimtime="00:02:18.62" />
                    <SPLIT distance="250" swimtime="00:02:48.68" />
                    <SPLIT distance="300" swimtime="00:03:21.29" />
                    <SPLIT distance="350" swimtime="00:03:50.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6906" number="1" />
                    <RELAYPOSITION athleteid="6945" number="2" />
                    <RELAYPOSITION athleteid="6934" number="3" />
                    <RELAYPOSITION athleteid="6919" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1399" points="521" swimtime="00:03:53.87" resultid="7072" heatid="10753" lane="3" entrytime="00:03:47.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.38" />
                    <SPLIT distance="100" swimtime="00:00:57.00" />
                    <SPLIT distance="150" swimtime="00:01:24.27" />
                    <SPLIT distance="200" swimtime="00:01:54.76" />
                    <SPLIT distance="250" swimtime="00:02:23.51" />
                    <SPLIT distance="300" swimtime="00:02:55.76" />
                    <SPLIT distance="350" swimtime="00:03:23.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6906" number="1" />
                    <RELAYPOSITION athleteid="6934" number="2" />
                    <RELAYPOSITION athleteid="6987" number="3" />
                    <RELAYPOSITION athleteid="6945" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1329" points="415" swimtime="00:04:37.17" resultid="7069" heatid="10697" lane="5" entrytime="00:04:27.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                    <SPLIT distance="100" swimtime="00:01:17.05" />
                    <SPLIT distance="150" swimtime="00:01:53.40" />
                    <SPLIT distance="200" swimtime="00:02:33.29" />
                    <SPLIT distance="250" swimtime="00:03:00.93" />
                    <SPLIT distance="300" swimtime="00:03:31.13" />
                    <SPLIT distance="350" swimtime="00:04:02.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6952" number="1" />
                    <RELAYPOSITION athleteid="6913" number="2" />
                    <RELAYPOSITION athleteid="6894" number="3" />
                    <RELAYPOSITION athleteid="6975" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1397" points="479" swimtime="00:04:00.57" resultid="7073" heatid="10752" lane="5" entrytime="00:04:01.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.96" />
                    <SPLIT distance="100" swimtime="00:00:53.28" />
                    <SPLIT distance="150" swimtime="00:01:21.43" />
                    <SPLIT distance="200" swimtime="00:01:52.30" />
                    <SPLIT distance="250" swimtime="00:02:24.06" />
                    <SPLIT distance="300" swimtime="00:02:58.76" />
                    <SPLIT distance="350" swimtime="00:03:28.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6894" number="1" />
                    <RELAYPOSITION athleteid="6952" number="2" />
                    <RELAYPOSITION athleteid="6975" number="3" />
                    <RELAYPOSITION athleteid="6913" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1323" points="306" swimtime="00:05:06.71" resultid="7070" heatid="10693" lane="6" entrytime="00:05:23.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.97" />
                    <SPLIT distance="100" swimtime="00:01:16.41" />
                    <SPLIT distance="150" swimtime="00:01:55.51" />
                    <SPLIT distance="200" swimtime="00:02:43.38" />
                    <SPLIT distance="250" swimtime="00:03:16.66" />
                    <SPLIT distance="300" swimtime="00:03:56.40" />
                    <SPLIT distance="350" swimtime="00:04:29.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7033" number="1" />
                    <RELAYPOSITION athleteid="7016" number="2" />
                    <RELAYPOSITION athleteid="7027" number="3" />
                    <RELAYPOSITION athleteid="7050" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1391" points="354" swimtime="00:04:25.99" resultid="7075" heatid="10748" lane="2" entrytime="00:04:25.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.19" />
                    <SPLIT distance="100" swimtime="00:01:05.88" />
                    <SPLIT distance="150" swimtime="00:01:38.49" />
                    <SPLIT distance="200" swimtime="00:02:13.45" />
                    <SPLIT distance="250" swimtime="00:02:46.47" />
                    <SPLIT distance="300" swimtime="00:03:24.33" />
                    <SPLIT distance="350" swimtime="00:03:54.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7033" number="1" />
                    <RELAYPOSITION athleteid="7016" number="2" />
                    <RELAYPOSITION athleteid="7039" number="3" />
                    <RELAYPOSITION athleteid="7027" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1325" points="326" swimtime="00:05:00.22" resultid="7071" heatid="10694" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                    <SPLIT distance="100" swimtime="00:01:09.21" />
                    <SPLIT distance="150" swimtime="00:01:49.94" />
                    <SPLIT distance="200" swimtime="00:02:34.29" />
                    <SPLIT distance="250" swimtime="00:03:10.89" />
                    <SPLIT distance="350" swimtime="00:04:25.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6900" number="1" />
                    <RELAYPOSITION athleteid="6981" number="2" />
                    <RELAYPOSITION athleteid="6925" number="3" />
                    <RELAYPOSITION athleteid="7061" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1393" points="395" swimtime="00:04:16.54" resultid="7074" heatid="10749" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.84" />
                    <SPLIT distance="100" swimtime="00:00:58.27" />
                    <SPLIT distance="150" swimtime="00:01:29.62" />
                    <SPLIT distance="200" swimtime="00:02:04.70" />
                    <SPLIT distance="250" swimtime="00:02:35.62" />
                    <SPLIT distance="300" swimtime="00:03:10.20" />
                    <SPLIT distance="350" swimtime="00:03:41.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6900" number="1" />
                    <RELAYPOSITION athleteid="6981" number="2" />
                    <RELAYPOSITION athleteid="6925" number="3" />
                    <RELAYPOSITION athleteid="7061" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1315" points="307" swimtime="00:05:40.27" resultid="7066" heatid="10689" lane="5" entrytime="00:05:14.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                    <SPLIT distance="150" swimtime="00:02:10.34" />
                    <SPLIT distance="200" swimtime="00:02:58.61" />
                    <SPLIT distance="250" swimtime="00:03:37.04" />
                    <SPLIT distance="300" swimtime="00:04:28.61" />
                    <SPLIT distance="350" swimtime="00:05:01.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7022" number="1" />
                    <RELAYPOSITION athleteid="7045" number="2" />
                    <RELAYPOSITION athleteid="7010" number="3" />
                    <RELAYPOSITION athleteid="7004" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1383" points="343" swimtime="00:04:56.93" resultid="7067" heatid="10744" lane="2" entrytime="00:04:39.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                    <SPLIT distance="100" swimtime="00:01:13.97" />
                    <SPLIT distance="150" swimtime="00:01:47.90" />
                    <SPLIT distance="200" swimtime="00:02:27.44" />
                    <SPLIT distance="250" swimtime="00:03:02.58" />
                    <SPLIT distance="300" swimtime="00:03:41.92" />
                    <SPLIT distance="350" swimtime="00:04:17.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7004" number="1" />
                    <RELAYPOSITION athleteid="7022" number="2" />
                    <RELAYPOSITION athleteid="7045" number="3" />
                    <RELAYPOSITION athleteid="7010" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1113" points="358" swimtime="00:05:05.96" resultid="7076" heatid="10510" lane="3" entrytime="00:04:52.99">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.50" />
                    <SPLIT distance="150" swimtime="00:02:00.89" />
                    <SPLIT distance="200" swimtime="00:02:43.81" />
                    <SPLIT distance="250" swimtime="00:03:15.78" />
                    <SPLIT distance="300" swimtime="00:03:52.85" />
                    <SPLIT distance="350" swimtime="00:04:25.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7010" number="1" />
                    <RELAYPOSITION athleteid="6981" number="2" />
                    <RELAYPOSITION athleteid="6900" number="3" />
                    <RELAYPOSITION athleteid="7004" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="X" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1111" points="332" swimtime="00:05:13.75" resultid="7077" heatid="10509" lane="3" entrytime="00:05:02.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.97" />
                    <SPLIT distance="100" swimtime="00:01:24.50" />
                    <SPLIT distance="150" swimtime="00:02:06.79" />
                    <SPLIT distance="200" swimtime="00:02:55.62" />
                    <SPLIT distance="250" swimtime="00:03:30.10" />
                    <SPLIT distance="300" swimtime="00:04:13.68" />
                    <SPLIT distance="350" swimtime="00:04:41.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7022" number="1" />
                    <RELAYPOSITION athleteid="7045" number="2" />
                    <RELAYPOSITION athleteid="7033" number="3" />
                    <RELAYPOSITION athleteid="7027" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="X" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1245" points="440" swimtime="00:04:45.71" resultid="7078" heatid="10630" lane="6" entrytime="00:04:46.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.48" />
                    <SPLIT distance="100" swimtime="00:01:22.41" />
                    <SPLIT distance="150" swimtime="00:01:58.82" />
                    <SPLIT distance="200" swimtime="00:02:38.80" />
                    <SPLIT distance="250" swimtime="00:03:05.72" />
                    <SPLIT distance="300" swimtime="00:03:35.25" />
                    <SPLIT distance="350" swimtime="00:04:07.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6993" number="1" />
                    <RELAYPOSITION athleteid="6913" number="2" />
                    <RELAYPOSITION athleteid="6894" number="3" />
                    <RELAYPOSITION athleteid="6940" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="15981" nation="BRA" region="PR" clubid="6556" swrid="93783" name="Quinto Nado" shortname="5º Nado">
          <ATHLETES>
            <ATHLETE firstname="Francisco" lastname="Silva Telles" birthdate="2011-07-19" gender="M" nation="BRA" license="377311" swrid="5603911" athleteid="6578" externalid="377311">
              <RESULTS>
                <RESULT eventid="1087" points="279" swimtime="00:03:11.90" resultid="6579" heatid="10488" lane="4" entrytime="00:03:19.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.71" />
                    <SPLIT distance="100" swimtime="00:01:32.97" />
                    <SPLIT distance="150" swimtime="00:02:25.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="322" swimtime="00:00:37.85" resultid="6580" heatid="10572" lane="8" entrytime="00:00:39.70" entrycourse="LCM" />
                <RESULT eventid="1155" points="307" swimtime="00:01:08.74" resultid="6581" heatid="10540" lane="5" entrytime="00:01:12.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="295" swimtime="00:01:25.44" resultid="6582" heatid="10593" lane="4" entrytime="00:01:29.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="297" swimtime="00:02:32.79" resultid="6583" heatid="10665" lane="2" entrytime="00:02:44.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                    <SPLIT distance="100" swimtime="00:01:12.74" />
                    <SPLIT distance="150" swimtime="00:01:53.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="326" swimtime="00:05:19.44" resultid="6584" heatid="10718" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                    <SPLIT distance="100" swimtime="00:01:15.40" />
                    <SPLIT distance="150" swimtime="00:01:56.38" />
                    <SPLIT distance="200" swimtime="00:02:37.85" />
                    <SPLIT distance="250" swimtime="00:03:19.33" />
                    <SPLIT distance="300" swimtime="00:04:00.98" />
                    <SPLIT distance="350" swimtime="00:04:42.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Kikuchi Fujii" birthdate="2007-01-04" gender="M" nation="BRA" license="297805" swrid="5603863" athleteid="6557" externalid="297805">
              <RESULTS>
                <RESULT eventid="1103" points="573" swimtime="00:00:26.81" resultid="6558" heatid="10508" lane="6" entrytime="00:00:26.45" entrycourse="LCM" />
                <RESULT eventid="1087" points="628" swimtime="00:02:26.51" resultid="6559" heatid="10492" lane="4" entrytime="00:02:22.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.93" />
                    <SPLIT distance="100" swimtime="00:01:09.81" />
                    <SPLIT distance="150" swimtime="00:01:48.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="575" swimtime="00:00:31.19" resultid="6560" heatid="10575" lane="2" entrytime="00:00:30.44" entrycourse="LCM" />
                <RESULT eventid="1219" points="586" swimtime="00:01:07.95" resultid="6561" heatid="10599" lane="7" entrytime="00:01:05.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="574" swimtime="00:02:17.10" resultid="6562" heatid="10652" lane="3" entrytime="00:02:15.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.64" />
                    <SPLIT distance="100" swimtime="00:01:05.00" />
                    <SPLIT distance="150" swimtime="00:01:45.40" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 9:27), Na volta dos 50m." eventid="1341" status="DSQ" swimtime="00:00:59.60" resultid="6563" heatid="10711" lane="6" entrytime="00:00:58.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Poletti Veiga" birthdate="2010-10-01" gender="F" nation="BRA" license="376951" swrid="5603895" athleteid="6564" externalid="376951">
              <RESULTS>
                <RESULT eventid="1063" points="408" swimtime="00:02:45.92" resultid="6565" heatid="10473" lane="9" entrytime="00:02:43.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                    <SPLIT distance="100" swimtime="00:01:20.55" />
                    <SPLIT distance="150" swimtime="00:02:03.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="547" swimtime="00:01:03.21" resultid="6566" heatid="10533" lane="1" entrytime="00:01:05.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="500" swimtime="00:00:29.73" resultid="6567" heatid="10607" lane="4" entrytime="00:00:29.82" entrycourse="LCM" />
                <RESULT eventid="1281" points="533" swimtime="00:02:18.36" resultid="6568" heatid="10660" lane="0" entrytime="00:02:19.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                    <SPLIT distance="100" swimtime="00:01:06.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="502" swimtime="00:04:56.16" resultid="6569" heatid="10716" lane="8" entrytime="00:05:02.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.71" />
                    <SPLIT distance="100" swimtime="00:01:11.57" />
                    <SPLIT distance="150" swimtime="00:01:50.10" />
                    <SPLIT distance="200" swimtime="00:02:28.45" />
                    <SPLIT distance="250" swimtime="00:03:06.24" />
                    <SPLIT distance="350" swimtime="00:04:20.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="412" swimtime="00:01:16.76" resultid="6570" heatid="10731" lane="8" entrytime="00:01:17.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Gomes" birthdate="2011-12-03" gender="F" nation="BRA" license="382051" swrid="5603846" athleteid="6585" externalid="382051">
              <RESULTS>
                <RESULT eventid="1179" points="103" swimtime="00:01:02.16" resultid="6586" heatid="10561" lane="8" />
                <RESULT eventid="1147" points="246" swimtime="00:01:22.42" resultid="6587" heatid="10524" lane="4" />
                <RESULT eventid="1227" points="270" swimtime="00:00:36.49" resultid="6588" heatid="10601" lane="5" entrytime="00:00:37.33" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Takemura Couto" birthdate="2010-02-08" gender="F" nation="BRA" license="376950" swrid="5603919" athleteid="6571" externalid="376950">
              <RESULTS>
                <RESULT eventid="1095" points="534" swimtime="00:00:30.11" resultid="6572" heatid="10498" lane="1" entrytime="00:00:31.88" entrycourse="LCM" />
                <RESULT eventid="1147" points="580" swimtime="00:01:02.00" resultid="6573" heatid="10533" lane="2" entrytime="00:01:05.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="586" swimtime="00:00:28.21" resultid="6574" heatid="10609" lane="9" entrytime="00:00:29.24" entrycourse="LCM" />
                <RESULT eventid="1281" points="491" swimtime="00:02:22.21" resultid="6575" heatid="10656" lane="8" entrytime="00:02:35.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                    <SPLIT distance="100" swimtime="00:01:06.67" />
                    <SPLIT distance="150" swimtime="00:01:44.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="380" swimtime="00:01:16.18" resultid="6576" heatid="10701" lane="8" entrytime="00:01:22.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="440" swimtime="00:01:15.08" resultid="6577" heatid="10730" lane="7" entrytime="00:01:19.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="11303" nation="BRA" region="PR" clubid="7279" swrid="93760" name="Associação De Talentos Da Natação" shortname="Atn/Curitiba">
          <ATHLETES>
            <ATHLETE firstname="Isaac" lastname="Zonta" birthdate="2012-11-14" gender="M" nation="BRA" license="414857" swrid="5755348" athleteid="7378" externalid="414857">
              <RESULTS>
                <RESULT eventid="1187" points="141" swimtime="00:00:49.79" resultid="7379" heatid="10570" lane="8" entrytime="00:00:51.89" entrycourse="LCM" />
                <RESULT eventid="1155" points="241" swimtime="00:01:14.50" resultid="7380" heatid="10539" lane="9" entrytime="00:01:16.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="246" swimtime="00:00:33.34" resultid="7381" heatid="10614" lane="3" entrytime="00:00:33.62" entrycourse="LCM" />
                <RESULT eventid="1219" points="130" swimtime="00:01:52.17" resultid="7382" heatid="10592" lane="9" entrytime="00:01:52.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Rosa Pech" birthdate="2010-10-26" gender="M" nation="BRA" license="413378" swrid="5755377" athleteid="7372" externalid="413378">
              <RESULTS>
                <RESULT eventid="1087" points="220" swimtime="00:03:27.62" resultid="7373" heatid="10488" lane="2" entrytime="00:03:26.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.00" />
                    <SPLIT distance="100" swimtime="00:01:40.78" />
                    <SPLIT distance="150" swimtime="00:02:34.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="266" swimtime="00:00:40.33" resultid="7374" heatid="10571" lane="6" entrytime="00:00:41.55" entrycourse="LCM" />
                <RESULT eventid="1155" points="250" swimtime="00:01:13.56" resultid="7375" heatid="10540" lane="6" entrytime="00:01:12.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="254" swimtime="00:00:32.98" resultid="7376" heatid="10613" lane="4" entrytime="00:00:35.73" entrycourse="LCM" />
                <RESULT eventid="1219" points="249" swimtime="00:01:30.31" resultid="7377" heatid="10593" lane="8" entrytime="00:01:33.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcos" lastname="Demchuk" birthdate="2011-06-15" gender="M" nation="BRA" license="388540" swrid="5602530" athleteid="7326" externalid="388540">
              <RESULTS>
                <RESULT eventid="1103" points="219" swimtime="00:00:36.93" resultid="7327" heatid="10502" lane="4" entrytime="00:00:38.55" entrycourse="LCM" />
                <RESULT eventid="1155" points="328" swimtime="00:01:07.25" resultid="7328" heatid="10543" lane="0" entrytime="00:01:07.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="314" swimtime="00:00:30.74" resultid="7329" heatid="10618" lane="4" entrytime="00:00:30.25" entrycourse="LCM" />
                <RESULT eventid="1289" points="269" swimtime="00:02:37.99" resultid="7330" heatid="10666" lane="8" entrytime="00:02:39.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                    <SPLIT distance="100" swimtime="00:01:11.47" />
                    <SPLIT distance="150" swimtime="00:01:54.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Arthur Ribeiro" birthdate="2010-02-05" gender="M" nation="BRA" license="408025" swrid="5723020" athleteid="7366" externalid="408025">
              <RESULTS>
                <RESULT eventid="1103" points="251" swimtime="00:00:35.30" resultid="7367" heatid="10503" lane="9" entrytime="00:00:37.30" entrycourse="LCM" />
                <RESULT eventid="1187" points="362" swimtime="00:00:36.38" resultid="7368" heatid="10574" lane="9" entrytime="00:00:35.49" entrycourse="LCM" />
                <RESULT eventid="1219" points="331" swimtime="00:01:22.20" resultid="7369" heatid="10595" lane="8" entrytime="00:01:23.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="244" swimtime="00:00:37.67" resultid="7370" heatid="10683" lane="1" />
                <RESULT eventid="1373" points="273" swimtime="00:01:19.49" resultid="7371" heatid="10735" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Zaleski Dallazem" birthdate="2009-05-16" gender="M" nation="BRA" license="344286" swrid="5600280" athleteid="7298" externalid="344286" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1087" points="432" swimtime="00:02:45.92" resultid="7299" heatid="10491" lane="2" entrytime="00:02:47.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                    <SPLIT distance="100" swimtime="00:01:19.54" />
                    <SPLIT distance="150" swimtime="00:02:02.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="469" swimtime="00:00:59.70" resultid="7300" heatid="10548" lane="5" entrytime="00:00:59.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="448" swimtime="00:01:14.33" resultid="7301" heatid="10597" lane="6" entrytime="00:01:14.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="420" swimtime="00:02:16.14" resultid="7302" heatid="10663" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.39" />
                    <SPLIT distance="100" swimtime="00:01:04.48" />
                    <SPLIT distance="150" swimtime="00:01:40.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Neves Vianna" birthdate="2007-12-30" gender="F" nation="BRA" license="391106" swrid="5600223" athleteid="7331" externalid="391106">
              <RESULTS>
                <RESULT eventid="1095" points="182" swimtime="00:00:43.07" resultid="7332" heatid="10495" lane="5" entrytime="00:00:44.61" entrycourse="LCM" />
                <RESULT eventid="1063" points="208" swimtime="00:03:27.73" resultid="7333" heatid="10470" lane="9" entrytime="00:03:20.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="246" swimtime="00:01:22.42" resultid="7334" heatid="10526" lane="7" entrytime="00:01:20.18" entrycourse="LCM" />
                <RESULT eventid="1297" points="240" swimtime="00:00:43.22" resultid="7335" heatid="10678" lane="1" entrytime="00:00:42.96" entrycourse="LCM" />
                <RESULT eventid="1281" points="217" swimtime="00:03:06.51" resultid="7336" heatid="10654" lane="2" entrytime="00:02:58.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.83" />
                    <SPLIT distance="100" swimtime="00:01:29.97" />
                    <SPLIT distance="150" swimtime="00:02:17.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="215" swimtime="00:01:35.26" resultid="7337" heatid="10727" lane="6" entrytime="00:01:32.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Santana Melosilva" birthdate="2008-08-18" gender="M" nation="BRA" license="421428" swrid="5638377" athleteid="7383" externalid="421428">
              <RESULTS>
                <RESULT eventid="1103" points="341" swimtime="00:00:31.87" resultid="7384" heatid="10504" lane="4" entrytime="00:00:33.19" entrycourse="LCM" />
                <RESULT eventid="1155" points="352" swimtime="00:01:05.71" resultid="7385" heatid="10542" lane="3" entrytime="00:01:09.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="364" swimtime="00:00:29.27" resultid="7386" heatid="10619" lane="5" entrytime="00:00:29.77" entrycourse="LCM" />
                <RESULT comment="SW 8.5 - Totalmente submerso durante o nado.  (Horário: 9:12)" eventid="1341" status="DSQ" swimtime="00:01:28.19" resultid="7387" heatid="10704" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Kerppers Kreia" birthdate="2006-12-01" gender="M" nation="BRA" license="366815" swrid="5600195" athleteid="7293" externalid="366815">
              <RESULTS>
                <RESULT eventid="1155" points="530" swimtime="00:00:57.31" resultid="7294" heatid="10550" lane="7" entrytime="00:00:57.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="478" swimtime="00:00:26.73" resultid="7295" heatid="10624" lane="2" entrytime="00:00:27.06" entrycourse="LCM" />
                <RESULT eventid="1289" points="510" swimtime="00:02:07.62" resultid="7296" heatid="10672" lane="3" entrytime="00:02:08.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.22" />
                    <SPLIT distance="100" swimtime="00:01:01.63" />
                    <SPLIT distance="150" swimtime="00:01:34.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="376" swimtime="00:01:08.51" resultid="7297" heatid="10708" lane="4" entrytime="00:01:07.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Camila" lastname="Duarte De Almeida" birthdate="2009-11-26" gender="F" nation="BRA" license="378819" swrid="5600152" athleteid="7315" externalid="378819">
              <RESULTS>
                <RESULT eventid="1095" points="383" swimtime="00:00:33.64" resultid="7316" heatid="10497" lane="5" entrytime="00:00:33.98" entrycourse="LCM" />
                <RESULT eventid="1179" points="324" swimtime="00:00:42.45" resultid="7317" heatid="10561" lane="3" />
                <RESULT eventid="1147" points="496" swimtime="00:01:05.30" resultid="7318" heatid="10532" lane="5" entrytime="00:01:05.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="501" swimtime="00:00:29.71" resultid="7319" heatid="10608" lane="7" entrytime="00:00:29.55" entrycourse="LCM" />
                <RESULT eventid="1297" points="404" swimtime="00:00:36.32" resultid="7320" heatid="10677" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Castellano Purkot" birthdate="2010-01-25" gender="M" nation="BRA" license="392484" swrid="5622268" athleteid="7338" externalid="392484">
              <RESULTS>
                <RESULT eventid="1187" points="249" swimtime="00:00:41.24" resultid="7339" heatid="10572" lane="0" entrytime="00:00:39.86" entrycourse="LCM" />
                <RESULT eventid="1155" points="337" swimtime="00:01:06.63" resultid="7340" heatid="10545" lane="2" entrytime="00:01:04.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="327" swimtime="00:00:30.35" resultid="7341" heatid="10620" lane="5" entrytime="00:00:29.36" entrycourse="LCM" />
                <RESULT eventid="1289" points="273" swimtime="00:02:37.21" resultid="7342" heatid="10663" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                    <SPLIT distance="100" swimtime="00:01:12.10" />
                    <SPLIT distance="150" swimtime="00:01:54.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabiana" lastname="Zaleski Dallazem" birthdate="2009-05-16" gender="F" nation="BRA" license="344287" swrid="5600279" athleteid="7280" externalid="344287">
              <RESULTS>
                <RESULT eventid="1063" points="512" swimtime="00:02:33.88" resultid="7281" heatid="10473" lane="3" entrytime="00:02:32.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                    <SPLIT distance="100" swimtime="00:01:14.55" />
                    <SPLIT distance="150" swimtime="00:01:53.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="518" swimtime="00:01:04.35" resultid="7282" heatid="10533" lane="5" entrytime="00:01:04.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="574" swimtime="00:00:32.31" resultid="7283" heatid="10680" lane="5" entrytime="00:00:32.05" entrycourse="LCM" />
                <RESULT comment="SW 6.5 - Não terminou a prova enquanto estava de costas.&#10;&#10;&#10;&#10;&#10;&#10;&#10;  (Horário: 16:22), Na volta dos 100m (Costas, Medley Individual)." eventid="1265" status="DSQ" swimtime="00:02:43.81" resultid="7284" heatid="10644" lane="2" entrytime="00:02:39.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                    <SPLIT distance="100" swimtime="00:01:15.39" />
                    <SPLIT distance="150" swimtime="00:02:06.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="562" swimtime="00:01:09.21" resultid="7285" heatid="10732" lane="5" entrytime="00:01:08.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Araujo Do Rego Barros" birthdate="2009-04-30" gender="M" nation="BRA" license="376325" swrid="5377739" athleteid="7303" externalid="376325">
              <RESULTS>
                <RESULT eventid="1103" points="379" swimtime="00:00:30.77" resultid="7304" heatid="10506" lane="1" entrytime="00:00:30.78" entrycourse="LCM" />
                <RESULT eventid="1171" points="338" swimtime="00:02:38.27" resultid="7305" heatid="10557" lane="1" entrytime="00:02:36.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                    <SPLIT distance="100" swimtime="00:01:11.97" />
                    <SPLIT distance="150" swimtime="00:01:54.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="408" swimtime="00:00:28.18" resultid="7306" heatid="10622" lane="8" entrytime="00:00:28.24" entrycourse="LCM" />
                <RESULT eventid="1273" points="328" swimtime="00:02:45.24" resultid="7307" heatid="10646" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.61" />
                    <SPLIT distance="100" swimtime="00:01:18.00" />
                    <SPLIT distance="150" swimtime="00:02:08.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="387" swimtime="00:01:07.82" resultid="7308" heatid="10708" lane="2" entrytime="00:01:08.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jhon" lastname="Caleb Dos Santos" birthdate="2010-03-02" gender="M" nation="BRA" license="359020" swrid="5588574" athleteid="7286" externalid="359020">
              <RESULTS>
                <RESULT eventid="1071" points="454" swimtime="00:02:25.57" resultid="7287" heatid="10475" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                    <SPLIT distance="100" swimtime="00:01:11.55" />
                    <SPLIT distance="150" swimtime="00:01:49.14" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 8.3 - Movimento alternado das pernas ou pés.  (Horário: 19:06)" eventid="1171" status="DSQ" swimtime="00:02:23.92" resultid="7288" heatid="10558" lane="0" entrytime="00:02:25.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                    <SPLIT distance="100" swimtime="00:01:05.21" />
                    <SPLIT distance="150" swimtime="00:01:42.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="445" swimtime="00:05:17.49" resultid="7289" heatid="10523" lane="9" entrytime="00:05:10.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                    <SPLIT distance="100" swimtime="00:01:09.50" />
                    <SPLIT distance="150" swimtime="00:01:50.79" />
                    <SPLIT distance="200" swimtime="00:02:31.50" />
                    <SPLIT distance="250" swimtime="00:03:20.02" />
                    <SPLIT distance="300" swimtime="00:04:07.49" />
                    <SPLIT distance="350" swimtime="00:04:43.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="538" swimtime="00:02:20.10" resultid="7290" heatid="10652" lane="1" entrytime="00:02:21.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.93" />
                    <SPLIT distance="100" swimtime="00:01:06.18" />
                    <SPLIT distance="150" swimtime="00:01:47.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="563" swimtime="00:00:59.88" resultid="7291" heatid="10711" lane="7" entrytime="00:00:59.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="558" swimtime="00:01:02.66" resultid="7292" heatid="10742" lane="0" entrytime="00:01:04.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Vinicius Zonta" birthdate="2012-11-14" gender="M" nation="BRA" license="399517" swrid="5652903" athleteid="7355" externalid="399517">
              <RESULTS>
                <RESULT eventid="1103" points="268" swimtime="00:00:34.52" resultid="7356" heatid="10503" lane="3" entrytime="00:00:35.34" entrycourse="LCM" />
                <RESULT eventid="1155" points="338" swimtime="00:01:06.57" resultid="7357" heatid="10543" lane="8" entrytime="00:01:07.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="334" swimtime="00:00:30.12" resultid="7358" heatid="10619" lane="9" entrytime="00:00:30.10" entrycourse="LCM" />
                <RESULT eventid="1289" points="267" swimtime="00:02:38.30" resultid="7359" heatid="10666" lane="0" entrytime="00:02:40.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="100" swimtime="00:01:14.06" />
                    <SPLIT distance="150" swimtime="00:01:56.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="194" swimtime="00:01:25.36" resultid="7360" heatid="10705" lane="6" entrytime="00:01:28.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Yuji Yamazato" birthdate="2008-10-01" gender="M" nation="BRA" license="392664" swrid="5622313" athleteid="7343" externalid="392664">
              <RESULTS>
                <RESULT eventid="1103" points="353" swimtime="00:00:31.50" resultid="7344" heatid="10506" lane="8" entrytime="00:00:30.83" entrycourse="LCM" />
                <RESULT eventid="1155" points="426" swimtime="00:01:01.66" resultid="7345" heatid="10547" lane="1" entrytime="00:01:01.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="429" swimtime="00:00:27.72" resultid="7346" heatid="10623" lane="7" entrytime="00:00:27.65" entrycourse="LCM" />
                <RESULT eventid="1305" points="361" swimtime="00:00:33.07" resultid="7347" heatid="10685" lane="2" entrytime="00:00:35.04" entrycourse="LCM" />
                <RESULT eventid="1373" points="336" swimtime="00:01:14.18" resultid="7348" heatid="10738" lane="5" entrytime="00:01:13.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yohanna" lastname="Vitoria Sena" birthdate="2012-01-20" gender="F" nation="BRA" license="406710" swrid="5717302" athleteid="7361" externalid="406710">
              <RESULTS>
                <RESULT eventid="1147" points="249" swimtime="00:01:22.17" resultid="7362" heatid="10525" lane="3" entrytime="00:01:22.06" entrycourse="LCM" />
                <RESULT eventid="1227" points="269" swimtime="00:00:36.56" resultid="7363" heatid="10602" lane="9" entrytime="00:00:37.03" entrycourse="LCM" />
                <RESULT eventid="1297" points="207" swimtime="00:00:45.36" resultid="7364" heatid="10678" lane="9" entrytime="00:00:45.87" entrycourse="LCM" />
                <RESULT eventid="1365" points="154" swimtime="00:01:46.46" resultid="7365" heatid="10726" lane="3" entrytime="00:01:50.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Fonseca Vendramin" birthdate="2008-09-28" gender="F" nation="BRA" license="393918" swrid="5622282" athleteid="7349" externalid="393918">
              <RESULTS>
                <RESULT eventid="1095" points="292" swimtime="00:00:36.81" resultid="7350" heatid="10497" lane="0" entrytime="00:00:36.31" entrycourse="LCM" />
                <RESULT eventid="1147" points="461" swimtime="00:01:06.90" resultid="7351" heatid="10530" lane="3" entrytime="00:01:08.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="416" swimtime="00:00:31.62" resultid="7352" heatid="10606" lane="3" entrytime="00:00:30.81" entrycourse="LCM" />
                <RESULT eventid="1297" points="419" swimtime="00:00:35.89" resultid="7353" heatid="10679" lane="4" entrytime="00:00:37.45" entrycourse="LCM" />
                <RESULT eventid="1365" points="350" swimtime="00:01:21.04" resultid="7354" heatid="10726" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Leal Kuss" birthdate="2012-10-20" gender="M" nation="BRA" license="385085" swrid="5588768" athleteid="7321" externalid="385085">
              <RESULTS>
                <RESULT eventid="1103" points="331" swimtime="00:00:32.19" resultid="7322" heatid="10504" lane="6" entrytime="00:00:33.43" entrycourse="LCM" />
                <RESULT eventid="1155" points="309" swimtime="00:01:08.57" resultid="7323" heatid="10541" lane="4" entrytime="00:01:10.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="312" swimtime="00:00:30.82" resultid="7324" heatid="10617" lane="0" entrytime="00:00:31.60" entrycourse="LCM" />
                <RESULT eventid="1341" points="239" swimtime="00:01:19.68" resultid="7325" heatid="10705" lane="4" entrytime="00:01:21.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Benetti Webber" birthdate="2008-12-10" gender="M" nation="BRA" license="421900" swrid="5820323" athleteid="7388" externalid="421900">
              <RESULTS>
                <RESULT eventid="1155" points="329" swimtime="00:01:07.20" resultid="7389" heatid="10543" lane="4" entrytime="00:01:06.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="379" swimtime="00:00:28.89" resultid="7390" heatid="10618" lane="2" entrytime="00:00:30.61" entrycourse="LCM" />
                <RESULT eventid="1289" points="252" swimtime="00:02:41.31" resultid="7391" heatid="10662" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                    <SPLIT distance="100" swimtime="00:01:11.92" />
                    <SPLIT distance="150" swimtime="00:01:56.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Muller" birthdate="2009-10-10" gender="F" nation="BRA" license="376952" swrid="5600221" athleteid="7309" externalid="376952">
              <RESULTS>
                <RESULT eventid="1079" points="450" swimtime="00:02:59.47" resultid="7310" heatid="10485" lane="1" entrytime="00:02:59.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.19" />
                    <SPLIT distance="100" swimtime="00:01:25.05" />
                    <SPLIT distance="150" swimtime="00:02:13.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="512" swimtime="00:00:36.44" resultid="7311" heatid="10565" lane="7" entrytime="00:00:36.39" entrycourse="LCM" />
                <RESULT eventid="1211" points="493" swimtime="00:01:21.16" resultid="7312" heatid="10589" lane="7" entrytime="00:01:19.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="444" swimtime="00:02:27.02" resultid="7313" heatid="10658" lane="2" entrytime="00:02:25.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.99" />
                    <SPLIT distance="100" swimtime="00:01:10.75" />
                    <SPLIT distance="150" swimtime="00:01:48.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="328" swimtime="00:01:22.81" resultid="7314" heatid="10726" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="ATN/CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1399" points="410" swimtime="00:04:13.20" resultid="7392" heatid="10753" lane="7" entrytime="00:03:56.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.72" />
                    <SPLIT distance="100" swimtime="00:00:57.53" />
                    <SPLIT distance="150" swimtime="00:01:26.44" />
                    <SPLIT distance="200" swimtime="00:01:58.99" />
                    <SPLIT distance="250" swimtime="00:02:29.91" />
                    <SPLIT distance="300" swimtime="00:03:05.85" />
                    <SPLIT distance="350" swimtime="00:03:36.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7293" number="1" />
                    <RELAYPOSITION athleteid="7343" number="2" />
                    <RELAYPOSITION athleteid="7388" number="3" />
                    <RELAYPOSITION athleteid="7383" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="ATN/CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT comment="SW 10.12 - Os pés perderam contato com a plataforma de partida antes que o colega de equipe anterior tocasse a borda.  (Horário: 13:11), Na volta dos 300m." eventid="1395" status="DSQ" swimtime="00:04:19.31" resultid="7393" heatid="10751" lane="5" entrytime="00:03:55.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.08" />
                    <SPLIT distance="100" swimtime="00:00:54.11" />
                    <SPLIT distance="150" swimtime="00:01:25.04" />
                    <SPLIT distance="200" swimtime="00:02:00.16" />
                    <SPLIT distance="250" swimtime="00:02:33.57" />
                    <SPLIT distance="350" swimtime="00:03:43.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7286" number="1" />
                    <RELAYPOSITION athleteid="7338" number="2" />
                    <RELAYPOSITION athleteid="7372" number="3" />
                    <RELAYPOSITION athleteid="7366" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="ATN/CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1393" points="312" swimtime="00:04:37.28" resultid="7394" heatid="10750" lane="7" entrytime="00:04:28.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                    <SPLIT distance="100" swimtime="00:01:09.39" />
                    <SPLIT distance="150" swimtime="00:01:39.70" />
                    <SPLIT distance="200" swimtime="00:02:15.15" />
                    <SPLIT distance="250" swimtime="00:02:49.34" />
                    <SPLIT distance="300" swimtime="00:03:28.33" />
                    <SPLIT distance="350" swimtime="00:04:00.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7326" number="1" />
                    <RELAYPOSITION athleteid="7355" number="2" />
                    <RELAYPOSITION athleteid="7378" number="3" />
                    <RELAYPOSITION athleteid="7321" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="X" name="ATN/CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1245" points="469" swimtime="00:04:39.77" resultid="7395" heatid="10630" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                    <SPLIT distance="100" swimtime="00:01:12.45" />
                    <SPLIT distance="150" swimtime="00:01:46.59" />
                    <SPLIT distance="200" swimtime="00:02:26.72" />
                    <SPLIT distance="250" swimtime="00:02:57.79" />
                    <SPLIT distance="300" swimtime="00:03:34.63" />
                    <SPLIT distance="350" swimtime="00:04:05.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="7280" number="1" />
                    <RELAYPOSITION athleteid="7298" number="2" />
                    <RELAYPOSITION athleteid="7303" number="3" />
                    <RELAYPOSITION athleteid="7315" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="1035" nation="BRA" region="PR" clubid="8760" swrid="93778" name="Fundação De Esportes De Campo Mourão" shortname="Fecam">
          <ATHLETES>
            <ATHLETE firstname="Julia" lastname="Gabrieli Oliveira" birthdate="2010-09-23" gender="F" nation="BRA" license="403428" swrid="5676288" athleteid="8798" externalid="403428">
              <RESULTS>
                <RESULT eventid="1147" points="274" swimtime="00:01:19.59" resultid="8799" heatid="10524" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="318" swimtime="00:00:34.58" resultid="8800" heatid="10601" lane="8" />
                <RESULT eventid="1297" points="217" swimtime="00:00:44.65" resultid="8801" heatid="10677" lane="8" />
                <RESULT eventid="1365" status="WDR" swimtime="00:00:00.00" resultid="8802" heatid="10726" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Ferreira Batista" birthdate="2012-03-29" gender="F" nation="BRA" license="385779" swrid="5532525" athleteid="8788" externalid="385779">
              <RESULTS>
                <RESULT eventid="1147" points="303" swimtime="00:01:16.93" resultid="8789" heatid="10524" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="316" swimtime="00:00:34.65" resultid="8790" heatid="10601" lane="9" />
                <RESULT eventid="1297" points="287" swimtime="00:00:40.68" resultid="8791" heatid="10677" lane="6" />
                <RESULT eventid="1365" points="246" swimtime="00:01:31.13" resultid="8792" heatid="10726" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kenzo" lastname="Kimura" birthdate="2010-04-23" gender="M" nation="BRA" license="403429" swrid="5676289" athleteid="8803" externalid="403429">
              <RESULTS>
                <RESULT eventid="1187" points="218" swimtime="00:00:43.10" resultid="8804" heatid="10567" lane="1" />
                <RESULT eventid="1155" points="276" swimtime="00:01:11.19" resultid="8805" heatid="10535" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="297" swimtime="00:00:31.34" resultid="8806" heatid="10610" lane="7" />
                <RESULT eventid="1289" points="219" swimtime="00:02:49.15" resultid="8807" heatid="10662" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                    <SPLIT distance="100" swimtime="00:01:14.63" />
                    <SPLIT distance="150" swimtime="00:02:02.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henry" lastname="Sadao Da Silva" birthdate="2012-10-02" gender="M" nation="BRA" license="413907" swrid="5755359" athleteid="8817" externalid="413907">
              <RESULTS>
                <RESULT eventid="1187" points="71" swimtime="00:01:02.50" resultid="8818" heatid="10568" lane="0" />
                <RESULT eventid="1155" points="143" swimtime="00:01:28.73" resultid="8819" heatid="10537" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="150" swimtime="00:00:39.33" resultid="8820" heatid="10612" lane="3" />
                <RESULT eventid="1373" points="106" swimtime="00:01:48.86" resultid="8821" heatid="10734" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Batinga Ponchielli" birthdate="2007-01-18" gender="M" nation="BRA" license="378461" swrid="5251143" athleteid="8776" externalid="378461">
              <RESULTS>
                <RESULT eventid="1155" points="282" swimtime="00:01:10.68" resultid="8777" heatid="10537" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="304" swimtime="00:00:31.09" resultid="8778" heatid="10613" lane="0" />
                <RESULT eventid="1305" points="288" swimtime="00:00:35.62" resultid="8779" heatid="10683" lane="8" />
                <RESULT eventid="1373" points="216" swimtime="00:01:25.94" resultid="8780" heatid="10735" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Capel Adelino" birthdate="2009-04-24" gender="M" nation="BRA" license="422154" swrid="5819267" athleteid="8822" externalid="422154">
              <RESULTS>
                <RESULT eventid="1155" points="190" swimtime="00:01:20.62" resultid="8823" heatid="10535" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="236" swimtime="00:00:33.80" resultid="8824" heatid="10610" lane="1" />
                <RESULT eventid="1305" points="152" swimtime="00:00:44.04" resultid="8825" heatid="10681" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Stipp Silva" birthdate="2009-12-02" gender="M" nation="BRA" license="378462" swrid="5603918" athleteid="8781" externalid="378462">
              <RESULTS>
                <RESULT eventid="1087" points="279" swimtime="00:03:11.89" resultid="8782" heatid="10487" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.74" />
                    <SPLIT distance="100" swimtime="00:01:31.22" />
                    <SPLIT distance="150" swimtime="00:02:24.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="436" swimtime="00:00:34.21" resultid="8783" heatid="10568" lane="8" />
                <RESULT eventid="1155" points="455" swimtime="00:01:00.30" resultid="8784" heatid="10546" lane="3" entrytime="00:01:02.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="482" swimtime="00:00:26.66" resultid="8785" heatid="10623" lane="4" entrytime="00:00:27.48" entrycourse="LCM" />
                <RESULT eventid="1219" points="343" swimtime="00:01:21.20" resultid="8786" heatid="10594" lane="7" entrytime="00:01:27.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="388" swimtime="00:02:19.80" resultid="8787" heatid="10667" lane="4" entrytime="00:02:27.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                    <SPLIT distance="100" swimtime="00:01:05.83" />
                    <SPLIT distance="150" swimtime="00:01:43.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Eduardo Schork Filho" birthdate="2012-12-28" gender="M" nation="BRA" license="413906" swrid="5755352" athleteid="8812" externalid="413906">
              <RESULTS>
                <RESULT eventid="1187" points="133" swimtime="00:00:50.75" resultid="8813" heatid="10567" lane="3" />
                <RESULT eventid="1155" points="159" swimtime="00:01:25.57" resultid="8814" heatid="10537" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="169" swimtime="00:00:37.80" resultid="8815" heatid="10612" lane="7" />
                <RESULT eventid="1219" points="142" swimtime="00:01:48.95" resultid="8816" heatid="10590" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Giroldo Santos" birthdate="2011-05-16" gender="M" nation="BRA" license="399602" swrid="5755354" athleteid="8808" externalid="399602">
              <RESULTS>
                <RESULT eventid="1155" points="217" swimtime="00:01:17.12" resultid="8809" heatid="10537" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="207" swimtime="00:00:35.30" resultid="8810" heatid="10611" lane="2" />
                <RESULT eventid="1373" points="155" swimtime="00:01:35.96" resultid="8811" heatid="10733" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Franca Rebollo" birthdate="2012-09-26" gender="M" nation="BRA" license="385780" swrid="5538081" athleteid="8761" externalid="385780">
              <RESULTS>
                <RESULT eventid="1155" points="160" swimtime="00:01:25.43" resultid="8762" heatid="10536" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="171" swimtime="00:00:37.65" resultid="8763" heatid="10613" lane="9" />
                <RESULT eventid="1305" points="127" swimtime="00:00:46.73" resultid="8764" heatid="10682" lane="2" />
                <RESULT eventid="1373" points="139" swimtime="00:01:39.43" resultid="8765" heatid="10734" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Samuel" lastname="Massuda Santos" birthdate="2012-06-09" gender="M" nation="BRA" license="392189" swrid="5603872" athleteid="8793" externalid="392189">
              <RESULTS>
                <RESULT eventid="1187" points="215" swimtime="00:00:43.31" resultid="8794" heatid="10568" lane="9" />
                <RESULT eventid="1305" points="217" swimtime="00:00:39.18" resultid="8795" heatid="10683" lane="7" />
                <RESULT eventid="1273" points="250" swimtime="00:03:00.77" resultid="8796" heatid="10645" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                    <SPLIT distance="100" swimtime="00:01:26.99" />
                    <SPLIT distance="150" swimtime="00:02:20.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="256" swimtime="00:01:21.18" resultid="8797" heatid="10735" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Keirrison" lastname="Leite Silva" birthdate="2011-08-02" gender="M" nation="BRA" license="392161" swrid="5603864" athleteid="8766" externalid="392161">
              <RESULTS>
                <RESULT eventid="1187" points="145" swimtime="00:00:49.31" resultid="8767" heatid="10568" lane="3" />
                <RESULT eventid="1155" points="153" swimtime="00:01:26.75" resultid="8768" heatid="10536" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="164" swimtime="00:00:38.18" resultid="8769" heatid="10612" lane="9" />
                <RESULT eventid="1305" points="90" swimtime="00:00:52.37" resultid="8770" heatid="10681" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique De Oliveira" birthdate="2009-07-28" gender="M" nation="BRA" license="414505" swrid="5755355" athleteid="8771" externalid="414505">
              <RESULTS>
                <RESULT eventid="1103" points="422" swimtime="00:00:29.68" resultid="8772" heatid="10501" lane="7" />
                <RESULT eventid="1155" points="402" swimtime="00:01:02.84" resultid="8773" heatid="10535" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="426" swimtime="00:00:27.77" resultid="8774" heatid="10612" lane="2" />
                <RESULT eventid="1289" points="305" swimtime="00:02:31.40" resultid="8775" heatid="10663" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.62" />
                    <SPLIT distance="100" swimtime="00:01:06.06" />
                    <SPLIT distance="150" swimtime="00:01:48.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" name="FECAM/PR &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1329" points="241" swimtime="00:05:32.16" resultid="8826" heatid="10697" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.44" />
                    <SPLIT distance="100" swimtime="00:01:45.90" />
                    <SPLIT distance="150" swimtime="00:02:23.03" />
                    <SPLIT distance="200" swimtime="00:03:08.34" />
                    <SPLIT distance="250" swimtime="00:03:39.79" />
                    <SPLIT distance="300" swimtime="00:04:22.66" />
                    <SPLIT distance="350" swimtime="00:04:54.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8822" number="1" />
                    <RELAYPOSITION athleteid="8781" number="2" />
                    <RELAYPOSITION athleteid="8771" number="3" />
                    <RELAYPOSITION athleteid="8803" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="SW 10.12 - Os pés perderam contato com a plataforma de partida antes que o colega de equipe anterior tocasse a borda.  (Horário: 13:17), Na volta dos 100m." eventid="1397" status="DSQ" swimtime="00:04:33.70" resultid="8828" heatid="10752" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.77" />
                    <SPLIT distance="100" swimtime="00:01:01.03" />
                    <SPLIT distance="150" swimtime="00:01:36.04" />
                    <SPLIT distance="200" swimtime="00:02:20.95" />
                    <SPLIT distance="250" swimtime="00:02:52.86" />
                    <SPLIT distance="300" swimtime="00:03:31.38" />
                    <SPLIT distance="350" swimtime="00:04:00.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8781" number="1" />
                    <RELAYPOSITION athleteid="8822" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="8803" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="8771" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="FECAM/PR &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1323" points="150" swimtime="00:06:28.87" resultid="8827" heatid="10693" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.77" />
                    <SPLIT distance="150" swimtime="00:02:31.12" />
                    <SPLIT distance="200" swimtime="00:03:30.00" />
                    <SPLIT distance="250" swimtime="00:04:09.17" />
                    <SPLIT distance="300" swimtime="00:05:00.39" />
                    <SPLIT distance="350" swimtime="00:05:40.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8761" number="1" />
                    <RELAYPOSITION athleteid="8812" number="2" />
                    <RELAYPOSITION athleteid="8793" number="3" />
                    <RELAYPOSITION athleteid="8817" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1391" points="167" swimtime="00:05:41.25" resultid="8829" heatid="10748" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                    <SPLIT distance="100" swimtime="00:01:14.26" />
                    <SPLIT distance="150" swimtime="00:01:55.41" />
                    <SPLIT distance="200" swimtime="00:02:41.30" />
                    <SPLIT distance="250" swimtime="00:03:23.73" />
                    <SPLIT distance="300" swimtime="00:04:11.93" />
                    <SPLIT distance="350" swimtime="00:04:52.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8793" number="1" />
                    <RELAYPOSITION athleteid="8761" number="2" />
                    <RELAYPOSITION athleteid="8812" number="3" />
                    <RELAYPOSITION athleteid="8817" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="16816" nation="BRA" region="SC" clubid="8865" swrid="94375" name="JURERê SPORTS CENTER" shortname="Jusc/Swimfloripa">
          <ATHLETES>
            <ATHLETE firstname="José" lastname="Roberto Vaz Guimarães Neto" birthdate="1996-11-14" gender="M" nation="BRA" license="109462" swrid="5206816" athleteid="8866" externalid="109462">
              <RESULTS>
                <RESULT eventid="1103" points="655" status="EXH" swimtime="00:00:25.64" resultid="8867" heatid="10508" lane="4" entrytime="00:00:24.66" entrycourse="LCM" />
                <RESULT eventid="1235" points="656" status="EXH" swimtime="00:00:24.06" resultid="8868" heatid="10628" lane="3" entrytime="00:00:23.54" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="1327" nation="BRA" region="SC" clubid="6589" swrid="93762" name="A. Jaraguaense De Ince. Nat. Competitiva" shortname="Ajinc">
          <ATHLETES>
            <ATHLETE firstname="Isabela" lastname="Hermenegildo" birthdate="2009-06-05" gender="F" nation="BRA" license="356022" swrid="5634667" athleteid="6642" externalid="356022">
              <RESULTS>
                <RESULT eventid="1063" points="379" status="EXH" swimtime="00:02:50.14" resultid="6643" heatid="10473" lane="8" entrytime="00:02:39.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="483" status="EXH" swimtime="00:01:05.89" resultid="6644" heatid="10533" lane="3" entrytime="00:01:04.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" status="WDR" swimtime="00:00:00.00" resultid="6645" heatid="10633" lane="4" entrytime="00:11:00.82" entrycourse="LCM" />
                <RESULT eventid="1227" status="WDR" swimtime="00:00:00.00" resultid="6646" heatid="10608" lane="0" entrytime="00:00:29.70" entrycourse="LCM" />
                <RESULT eventid="1265" status="WDR" swimtime="00:00:00.00" resultid="6647" heatid="10642" lane="1" entrytime="00:02:51.44" entrycourse="LCM" />
                <RESULT eventid="1349" status="WDR" swimtime="00:00:00.00" resultid="6648" heatid="10715" lane="5" entrytime="00:05:05.35" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariana" lastname="Maestri Lima" birthdate="2011-06-06" gender="F" nation="BRA" license="394879" athleteid="6782" externalid="394879">
              <RESULTS>
                <RESULT eventid="1079" points="312" status="EXH" swimtime="00:03:22.60" resultid="6783" heatid="10483" lane="0" entrytime="00:03:17.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.86" />
                    <SPLIT distance="100" swimtime="00:01:34.24" />
                    <SPLIT distance="150" swimtime="00:02:28.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="380" status="EXH" swimtime="00:01:11.36" resultid="6784" heatid="10529" lane="8" entrytime="00:01:12.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="306" status="EXH" swimtime="00:01:35.11" resultid="6785" heatid="10585" lane="0" entrytime="00:01:33.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="364" status="EXH" swimtime="00:02:37.11" resultid="6786" heatid="10655" lane="6" entrytime="00:02:38.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                    <SPLIT distance="100" swimtime="00:01:12.75" />
                    <SPLIT distance="150" swimtime="00:01:54.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="340" status="EXH" swimtime="00:05:37.09" resultid="6787" heatid="10713" lane="2" entrytime="00:05:35.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                    <SPLIT distance="100" swimtime="00:01:17.00" />
                    <SPLIT distance="150" swimtime="00:01:59.26" />
                    <SPLIT distance="200" swimtime="00:02:42.99" />
                    <SPLIT distance="250" swimtime="00:03:26.82" />
                    <SPLIT distance="300" swimtime="00:04:10.79" />
                    <SPLIT distance="350" swimtime="00:04:53.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="322" status="EXH" swimtime="00:01:23.34" resultid="6788" heatid="10729" lane="6" entrytime="00:01:22.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kiara" lastname="Barauna Sagaz" birthdate="2007-06-13" gender="F" nation="BRA" license="331781" swrid="5634531" athleteid="6621" externalid="331781">
              <RESULTS>
                <RESULT eventid="1063" points="408" status="EXH" swimtime="00:02:45.97" resultid="6622" heatid="10472" lane="3" entrytime="00:02:45.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                    <SPLIT distance="100" swimtime="00:01:19.11" />
                    <SPLIT distance="150" swimtime="00:02:02.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="488" status="EXH" swimtime="00:01:05.64" resultid="6623" heatid="10524" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="499" status="EXH" swimtime="00:00:29.76" resultid="6624" heatid="10608" lane="6" entrytime="00:00:29.33" entrycourse="LCM" />
                <RESULT eventid="1211" points="381" status="EXH" swimtime="00:01:28.42" resultid="6625" heatid="10586" lane="3" entrytime="00:01:27.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="396" status="EXH" swimtime="00:02:51.69" resultid="6626" heatid="10642" lane="4" entrytime="00:02:49.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.60" />
                    <SPLIT distance="100" swimtime="00:01:20.03" />
                    <SPLIT distance="150" swimtime="00:02:10.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="418" status="EXH" swimtime="00:01:16.35" resultid="6627" heatid="10731" lane="4" entrytime="00:01:14.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Possamai" birthdate="2010-07-12" gender="F" nation="BRA" license="358444" swrid="5588865" athleteid="6663" externalid="358444">
              <RESULTS>
                <RESULT eventid="1079" points="402" status="EXH" swimtime="00:03:06.35" resultid="6664" heatid="10484" lane="4" entrytime="00:03:03.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.03" />
                    <SPLIT distance="100" swimtime="00:01:29.81" />
                    <SPLIT distance="150" swimtime="00:02:19.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="388" status="EXH" swimtime="00:06:02.34" resultid="6665" heatid="10520" lane="2" entrytime="00:05:49.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                    <SPLIT distance="100" swimtime="00:01:23.59" />
                    <SPLIT distance="150" swimtime="00:02:10.90" />
                    <SPLIT distance="200" swimtime="00:02:56.00" />
                    <SPLIT distance="250" swimtime="00:03:45.56" />
                    <SPLIT distance="300" swimtime="00:04:37.67" />
                    <SPLIT distance="350" swimtime="00:05:20.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="394" status="EXH" swimtime="00:01:27.47" resultid="6666" heatid="10587" lane="8" entrytime="00:01:26.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="441" status="EXH" swimtime="00:02:45.60" resultid="6667" heatid="10643" lane="4" entrytime="00:02:42.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="100" swimtime="00:01:18.33" />
                    <SPLIT distance="150" swimtime="00:02:06.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="332" status="EXH" swimtime="00:01:19.62" resultid="6668" heatid="10701" lane="6" entrytime="00:01:17.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="395" status="EXH" swimtime="00:01:17.82" resultid="6669" heatid="10725" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Erick" lastname="Lima" birthdate="2008-09-02" gender="M" nation="BRA" license="341465" swrid="5634688" athleteid="6628" externalid="341465">
              <RESULTS>
                <RESULT eventid="1123" points="491" status="EXH" swimtime="00:09:33.00" resultid="6629" heatid="10513" lane="0" entrytime="00:09:13.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                    <SPLIT distance="100" swimtime="00:01:05.63" />
                    <SPLIT distance="150" swimtime="00:01:40.75" />
                    <SPLIT distance="200" swimtime="00:02:15.77" />
                    <SPLIT distance="250" swimtime="00:02:51.41" />
                    <SPLIT distance="300" swimtime="00:03:27.41" />
                    <SPLIT distance="350" swimtime="00:04:03.83" />
                    <SPLIT distance="400" swimtime="00:04:40.63" />
                    <SPLIT distance="450" swimtime="00:05:17.21" />
                    <SPLIT distance="500" swimtime="00:05:54.41" />
                    <SPLIT distance="550" swimtime="00:06:31.13" />
                    <SPLIT distance="600" swimtime="00:07:07.99" />
                    <SPLIT distance="650" swimtime="00:07:44.67" />
                    <SPLIT distance="700" swimtime="00:08:21.09" />
                    <SPLIT distance="750" swimtime="00:08:57.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="475" status="EXH" swimtime="00:02:23.40" resultid="6630" heatid="10479" lane="7" entrytime="00:02:26.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                    <SPLIT distance="150" swimtime="00:01:47.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="449" status="EXH" swimtime="00:05:16.49" resultid="6631" heatid="10522" lane="5" entrytime="00:05:13.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="100" swimtime="00:01:12.76" />
                    <SPLIT distance="150" swimtime="00:01:52.66" />
                    <SPLIT distance="200" swimtime="00:02:31.22" />
                    <SPLIT distance="250" swimtime="00:03:20.43" />
                    <SPLIT distance="300" swimtime="00:04:09.18" />
                    <SPLIT distance="350" swimtime="00:04:43.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="502" status="EXH" swimtime="00:18:14.91" resultid="6632" heatid="10635" lane="3" entrytime="00:17:24.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                    <SPLIT distance="100" swimtime="00:01:08.34" />
                    <SPLIT distance="150" swimtime="00:01:43.62" />
                    <SPLIT distance="200" swimtime="00:02:19.25" />
                    <SPLIT distance="250" swimtime="00:02:54.73" />
                    <SPLIT distance="300" swimtime="00:03:30.84" />
                    <SPLIT distance="350" swimtime="00:04:07.16" />
                    <SPLIT distance="400" swimtime="00:04:44.23" />
                    <SPLIT distance="450" swimtime="00:05:20.78" />
                    <SPLIT distance="500" swimtime="00:05:57.99" />
                    <SPLIT distance="550" swimtime="00:06:34.79" />
                    <SPLIT distance="600" swimtime="00:07:12.08" />
                    <SPLIT distance="650" swimtime="00:07:49.41" />
                    <SPLIT distance="700" swimtime="00:08:27.03" />
                    <SPLIT distance="750" swimtime="00:09:04.28" />
                    <SPLIT distance="800" swimtime="00:09:42.11" />
                    <SPLIT distance="850" swimtime="00:10:19.44" />
                    <SPLIT distance="900" swimtime="00:10:57.28" />
                    <SPLIT distance="950" swimtime="00:11:34.68" />
                    <SPLIT distance="1000" swimtime="00:12:12.16" />
                    <SPLIT distance="1050" swimtime="00:12:49.53" />
                    <SPLIT distance="1100" swimtime="00:13:26.73" />
                    <SPLIT distance="1150" swimtime="00:14:03.13" />
                    <SPLIT distance="1200" swimtime="00:14:39.78" />
                    <SPLIT distance="1250" swimtime="00:15:16.28" />
                    <SPLIT distance="1300" swimtime="00:15:52.84" />
                    <SPLIT distance="1350" swimtime="00:16:29.00" />
                    <SPLIT distance="1400" swimtime="00:17:05.31" />
                    <SPLIT distance="1450" swimtime="00:17:40.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="482" status="EXH" swimtime="00:02:10.06" resultid="6633" heatid="10673" lane="1" entrytime="00:02:06.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.86" />
                    <SPLIT distance="100" swimtime="00:01:03.02" />
                    <SPLIT distance="150" swimtime="00:01:37.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="538" status="EXH" swimtime="00:04:30.49" resultid="6634" heatid="10724" lane="9" entrytime="00:04:27.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                    <SPLIT distance="100" swimtime="00:01:03.93" />
                    <SPLIT distance="150" swimtime="00:01:37.55" />
                    <SPLIT distance="200" swimtime="00:02:11.65" />
                    <SPLIT distance="250" swimtime="00:02:45.76" />
                    <SPLIT distance="300" swimtime="00:03:20.77" />
                    <SPLIT distance="350" swimtime="00:03:55.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emily" lastname="Dos Santos Jahn" birthdate="2012-10-22" gender="F" nation="BRA" license="405087" athleteid="6796" externalid="405087">
              <RESULTS>
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 10:07), Na volta dos 100m." eventid="1079" status="DSQ" swimtime="00:03:32.38" resultid="6797" heatid="10482" lane="6" entrytime="00:03:28.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.46" />
                    <SPLIT distance="100" swimtime="00:01:41.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="311" status="EXH" swimtime="00:00:43.01" resultid="6798" heatid="10562" lane="5" entrytime="00:00:43.45" entrycourse="LCM" />
                <RESULT eventid="1211" points="295" status="EXH" swimtime="00:01:36.27" resultid="6799" heatid="10585" lane="8" entrytime="00:01:33.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="295" status="EXH" swimtime="00:03:09.32" resultid="6800" heatid="10640" lane="4" entrytime="00:03:09.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.45" />
                    <SPLIT distance="150" swimtime="00:02:26.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="274" status="EXH" swimtime="00:02:52.70" resultid="6801" heatid="10653" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.78" />
                    <SPLIT distance="100" swimtime="00:01:25.06" />
                    <SPLIT distance="150" swimtime="00:02:09.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="272" status="EXH" swimtime="00:01:28.13" resultid="6802" heatid="10728" lane="8" entrytime="00:01:29.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucca" lastname="Pereira Ferronatto" birthdate="2011-03-31" gender="M" nation="BRA" license="367950" swrid="5627328" athleteid="6705" externalid="367950">
              <RESULTS>
                <RESULT eventid="1071" points="396" status="EXH" swimtime="00:02:32.39" resultid="6706" heatid="10478" lane="6" entrytime="00:02:29.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                    <SPLIT distance="100" swimtime="00:01:12.08" />
                    <SPLIT distance="150" swimtime="00:01:51.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="443" status="EXH" swimtime="00:01:00.83" resultid="6707" heatid="10548" lane="3" entrytime="00:01:00.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="408" status="EXH" swimtime="00:00:28.18" resultid="6708" heatid="10624" lane="9" entrytime="00:00:27.47" entrycourse="LCM" />
                <RESULT eventid="1273" points="401" status="EXH" swimtime="00:02:34.47" resultid="6709" heatid="10650" lane="2" entrytime="00:02:32.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                    <SPLIT distance="100" swimtime="00:01:12.06" />
                    <SPLIT distance="150" swimtime="00:02:00.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="405" status="EXH" swimtime="00:02:17.75" resultid="6710" heatid="10662" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.19" />
                    <SPLIT distance="100" swimtime="00:01:06.73" />
                    <SPLIT distance="150" swimtime="00:01:42.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="422" status="EXH" swimtime="00:01:08.77" resultid="6711" heatid="10740" lane="6" entrytime="00:01:07.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduarda" lastname="Possamai Da Silva" birthdate="2011-03-26" gender="F" nation="BRA" license="367939" swrid="5627342" athleteid="6684" externalid="367939">
              <RESULTS>
                <RESULT eventid="1115" points="376" status="EXH" swimtime="00:21:14.19" resultid="6685" heatid="10512" lane="6" entrytime="00:20:57.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                    <SPLIT distance="100" swimtime="00:01:18.11" />
                    <SPLIT distance="150" swimtime="00:01:59.47" />
                    <SPLIT distance="200" swimtime="00:02:41.39" />
                    <SPLIT distance="250" swimtime="00:03:23.56" />
                    <SPLIT distance="300" swimtime="00:04:06.27" />
                    <SPLIT distance="350" swimtime="00:04:48.60" />
                    <SPLIT distance="400" swimtime="00:05:31.15" />
                    <SPLIT distance="450" swimtime="00:06:13.33" />
                    <SPLIT distance="500" swimtime="00:06:56.09" />
                    <SPLIT distance="550" swimtime="00:07:38.70" />
                    <SPLIT distance="600" swimtime="00:08:21.24" />
                    <SPLIT distance="650" swimtime="00:09:04.32" />
                    <SPLIT distance="700" swimtime="00:09:47.35" />
                    <SPLIT distance="750" swimtime="00:10:30.51" />
                    <SPLIT distance="800" swimtime="00:11:14.03" />
                    <SPLIT distance="850" swimtime="00:11:56.71" />
                    <SPLIT distance="900" swimtime="00:12:39.83" />
                    <SPLIT distance="950" swimtime="00:13:23.20" />
                    <SPLIT distance="1000" swimtime="00:14:06.27" />
                    <SPLIT distance="1050" swimtime="00:14:49.40" />
                    <SPLIT distance="1100" swimtime="00:15:32.74" />
                    <SPLIT distance="1150" swimtime="00:16:15.96" />
                    <SPLIT distance="1200" swimtime="00:16:59.15" />
                    <SPLIT distance="1250" swimtime="00:17:41.71" />
                    <SPLIT distance="1300" swimtime="00:18:24.92" />
                    <SPLIT distance="1350" swimtime="00:19:07.55" />
                    <SPLIT distance="1400" swimtime="00:19:50.54" />
                    <SPLIT distance="1450" swimtime="00:20:33.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="393" status="EXH" swimtime="00:03:07.71" resultid="6686" heatid="10483" lane="5" entrytime="00:03:12.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                    <SPLIT distance="100" swimtime="00:01:29.85" />
                    <SPLIT distance="150" swimtime="00:02:20.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="381" status="EXH" swimtime="00:11:08.67" resultid="6687" heatid="10633" lane="6" entrytime="00:11:28.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                    <SPLIT distance="100" swimtime="00:01:12.37" />
                    <SPLIT distance="150" swimtime="00:01:53.20" />
                    <SPLIT distance="200" swimtime="00:02:35.58" />
                    <SPLIT distance="250" swimtime="00:03:17.80" />
                    <SPLIT distance="300" swimtime="00:04:01.60" />
                    <SPLIT distance="350" swimtime="00:04:44.27" />
                    <SPLIT distance="400" swimtime="00:05:27.44" />
                    <SPLIT distance="450" swimtime="00:06:10.60" />
                    <SPLIT distance="500" swimtime="00:06:54.06" />
                    <SPLIT distance="550" swimtime="00:07:37.38" />
                    <SPLIT distance="600" swimtime="00:08:20.48" />
                    <SPLIT distance="650" swimtime="00:09:03.16" />
                    <SPLIT distance="700" swimtime="00:09:46.66" />
                    <SPLIT distance="750" swimtime="00:10:28.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="423" status="EXH" swimtime="00:01:25.43" resultid="6688" heatid="10586" lane="5" entrytime="00:01:27.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="393" status="EXH" swimtime="00:02:33.09" resultid="6689" heatid="10655" lane="5" entrytime="00:02:37.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:11.23" />
                    <SPLIT distance="150" swimtime="00:01:52.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="387" status="EXH" swimtime="00:05:22.95" resultid="6690" heatid="10713" lane="6" entrytime="00:05:34.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                    <SPLIT distance="100" swimtime="00:01:13.44" />
                    <SPLIT distance="150" swimtime="00:01:54.09" />
                    <SPLIT distance="200" swimtime="00:02:35.26" />
                    <SPLIT distance="250" swimtime="00:03:17.14" />
                    <SPLIT distance="300" swimtime="00:04:00.14" />
                    <SPLIT distance="350" swimtime="00:04:41.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lara" lastname="Jacob Goncalves" birthdate="2011-02-26" gender="F" nation="BRA" license="405088" athleteid="6803" externalid="405088">
              <RESULTS>
                <RESULT eventid="1079" points="403" status="EXH" swimtime="00:03:06.11" resultid="6804" heatid="10484" lane="6" entrytime="00:03:05.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.86" />
                    <SPLIT distance="100" swimtime="00:01:29.90" />
                    <SPLIT distance="150" swimtime="00:02:19.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="405" status="EXH" swimtime="00:00:39.41" resultid="6805" heatid="10564" lane="1" entrytime="00:00:38.95" entrycourse="LCM" />
                <RESULT eventid="1131" points="275" status="EXH" swimtime="00:06:46.46" resultid="6806" heatid="10518" lane="4" entrytime="00:06:32.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.07" />
                    <SPLIT distance="100" swimtime="00:01:45.17" />
                    <SPLIT distance="150" swimtime="00:02:39.52" />
                    <SPLIT distance="200" swimtime="00:03:33.23" />
                    <SPLIT distance="250" swimtime="00:04:23.35" />
                    <SPLIT distance="300" swimtime="00:05:13.09" />
                    <SPLIT distance="350" swimtime="00:06:00.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="417" status="EXH" swimtime="00:01:25.79" resultid="6807" heatid="10587" lane="3" entrytime="00:01:24.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="310" status="EXH" swimtime="00:03:06.16" resultid="6808" heatid="10641" lane="7" entrytime="00:03:01.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.41" />
                    <SPLIT distance="100" swimtime="00:01:33.65" />
                    <SPLIT distance="150" swimtime="00:02:22.66" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 8.3 - Movimento alternado das pernas ou pés.  (Horário: 9:02)" eventid="1333" status="DSQ" swimtime="00:01:38.77" resultid="6809" heatid="10700" lane="7" entrytime="00:01:29.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Magalhães Brando" birthdate="2012-01-27" gender="M" nation="BRA" license="422941" athleteid="6810" externalid="422941">
              <RESULTS>
                <RESULT eventid="1071" points="188" status="EXH" swimtime="00:03:15.33" resultid="6811" heatid="10475" lane="5" entrytime="00:03:15.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.00" />
                    <SPLIT distance="100" swimtime="00:01:37.50" />
                    <SPLIT distance="150" swimtime="00:02:26.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="264" status="EXH" swimtime="00:01:12.30" resultid="6812" heatid="10539" lane="5" entrytime="00:01:14.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="289" status="EXH" swimtime="00:00:31.60" resultid="6813" heatid="10612" lane="6" />
                <RESULT eventid="1219" points="167" status="EXH" swimtime="00:01:43.15" resultid="6814" heatid="10592" lane="1" entrytime="00:01:42.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="246" status="EXH" swimtime="00:02:42.78" resultid="6815" heatid="10665" lane="8" entrytime="00:02:47.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                    <SPLIT distance="100" swimtime="00:01:20.64" />
                    <SPLIT distance="150" swimtime="00:02:03.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="219" status="EXH" swimtime="00:01:25.53" resultid="6816" heatid="10735" lane="4" entrytime="00:01:26.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cecília" lastname="CORRêA DE LIMA" birthdate="2012-05-08" gender="F" nation="BRA" license="369470" swrid="5748647" athleteid="6712" externalid="369470">
              <RESULTS>
                <RESULT eventid="1147" points="502" status="EXH" swimtime="00:01:05.05" resultid="6713" heatid="10534" lane="9" entrytime="00:01:04.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="387" status="EXH" swimtime="00:06:02.61" resultid="6714" heatid="10520" lane="1" entrytime="00:05:57.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.97" />
                    <SPLIT distance="100" swimtime="00:01:22.34" />
                    <SPLIT distance="150" swimtime="00:02:10.57" />
                    <SPLIT distance="200" swimtime="00:02:57.35" />
                    <SPLIT distance="250" swimtime="00:03:50.34" />
                    <SPLIT distance="300" swimtime="00:04:42.32" />
                    <SPLIT distance="350" swimtime="00:05:23.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="462" status="EXH" swimtime="00:10:26.80" resultid="6715" heatid="10632" lane="1" entrytime="00:10:38.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                    <SPLIT distance="100" swimtime="00:01:12.66" />
                    <SPLIT distance="150" swimtime="00:01:51.27" />
                    <SPLIT distance="200" swimtime="00:02:30.84" />
                    <SPLIT distance="250" swimtime="00:03:10.58" />
                    <SPLIT distance="300" swimtime="00:03:50.68" />
                    <SPLIT distance="350" swimtime="00:04:30.61" />
                    <SPLIT distance="400" swimtime="00:05:10.32" />
                    <SPLIT distance="450" swimtime="00:05:50.14" />
                    <SPLIT distance="500" swimtime="00:06:30.41" />
                    <SPLIT distance="550" swimtime="00:07:10.49" />
                    <SPLIT distance="600" swimtime="00:07:50.80" />
                    <SPLIT distance="650" swimtime="00:08:30.70" />
                    <SPLIT distance="700" swimtime="00:09:09.83" />
                    <SPLIT distance="750" swimtime="00:09:48.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="429" status="EXH" swimtime="00:02:47.14" resultid="6716" heatid="10643" lane="0" entrytime="00:02:47.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                    <SPLIT distance="100" swimtime="00:01:18.91" />
                    <SPLIT distance="150" swimtime="00:02:09.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="488" status="EXH" swimtime="00:02:22.48" resultid="6717" heatid="10659" lane="0" entrytime="00:02:23.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.78" />
                    <SPLIT distance="100" swimtime="00:01:08.24" />
                    <SPLIT distance="150" swimtime="00:01:45.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="478" status="EXH" swimtime="00:05:00.97" resultid="6718" heatid="10716" lane="9" entrytime="00:05:03.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="100" swimtime="00:01:11.73" />
                    <SPLIT distance="150" swimtime="00:01:49.84" />
                    <SPLIT distance="200" swimtime="00:02:28.44" />
                    <SPLIT distance="250" swimtime="00:03:06.83" />
                    <SPLIT distance="300" swimtime="00:03:45.00" />
                    <SPLIT distance="350" swimtime="00:04:23.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Fructuozo De Freitas" birthdate="2011-03-03" gender="M" nation="BRA" license="367946" swrid="5627252" athleteid="6691" externalid="367946">
              <RESULTS>
                <RESULT eventid="1123" points="394" status="EXH" swimtime="00:10:16.53" resultid="6692" heatid="10514" lane="0" entrytime="00:09:59.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                    <SPLIT distance="100" swimtime="00:01:10.16" />
                    <SPLIT distance="150" swimtime="00:01:47.47" />
                    <SPLIT distance="200" swimtime="00:02:25.53" />
                    <SPLIT distance="250" swimtime="00:03:05.08" />
                    <SPLIT distance="300" swimtime="00:03:44.34" />
                    <SPLIT distance="350" swimtime="00:04:23.76" />
                    <SPLIT distance="400" swimtime="00:05:02.99" />
                    <SPLIT distance="450" swimtime="00:05:43.32" />
                    <SPLIT distance="500" swimtime="00:06:22.05" />
                    <SPLIT distance="550" swimtime="00:07:02.49" />
                    <SPLIT distance="600" swimtime="00:07:42.14" />
                    <SPLIT distance="650" swimtime="00:08:22.01" />
                    <SPLIT distance="700" swimtime="00:09:00.89" />
                    <SPLIT distance="750" swimtime="00:09:40.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="415" status="EXH" swimtime="00:02:27.87" resultid="6693" heatid="10558" lane="9" entrytime="00:02:25.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                    <SPLIT distance="100" swimtime="00:01:08.62" />
                    <SPLIT distance="150" swimtime="00:01:48.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="394" status="EXH" swimtime="00:19:46.73" resultid="6694" heatid="10636" lane="9" entrytime="00:19:36.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.99" />
                    <SPLIT distance="100" swimtime="00:01:11.55" />
                    <SPLIT distance="150" swimtime="00:01:50.13" />
                    <SPLIT distance="200" swimtime="00:02:28.30" />
                    <SPLIT distance="250" swimtime="00:03:06.29" />
                    <SPLIT distance="300" swimtime="00:03:45.96" />
                    <SPLIT distance="350" swimtime="00:04:24.85" />
                    <SPLIT distance="400" swimtime="00:05:03.95" />
                    <SPLIT distance="450" swimtime="00:05:43.09" />
                    <SPLIT distance="500" swimtime="00:06:22.19" />
                    <SPLIT distance="550" swimtime="00:07:01.62" />
                    <SPLIT distance="600" swimtime="00:07:41.58" />
                    <SPLIT distance="650" swimtime="00:08:20.74" />
                    <SPLIT distance="700" swimtime="00:09:00.64" />
                    <SPLIT distance="750" swimtime="00:09:39.68" />
                    <SPLIT distance="800" swimtime="00:10:20.04" />
                    <SPLIT distance="850" swimtime="00:10:59.56" />
                    <SPLIT distance="900" swimtime="00:11:40.47" />
                    <SPLIT distance="950" swimtime="00:12:20.18" />
                    <SPLIT distance="1000" swimtime="00:13:01.05" />
                    <SPLIT distance="1050" swimtime="00:13:41.15" />
                    <SPLIT distance="1100" swimtime="00:14:22.15" />
                    <SPLIT distance="1150" swimtime="00:15:02.58" />
                    <SPLIT distance="1200" swimtime="00:15:43.56" />
                    <SPLIT distance="1250" swimtime="00:16:24.29" />
                    <SPLIT distance="1300" swimtime="00:17:05.27" />
                    <SPLIT distance="1350" swimtime="00:17:45.57" />
                    <SPLIT distance="1400" swimtime="00:18:26.51" />
                    <SPLIT distance="1450" swimtime="00:19:06.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="343" status="EXH" swimtime="00:02:42.85" resultid="6695" heatid="10649" lane="3" entrytime="00:02:38.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                    <SPLIT distance="100" swimtime="00:01:16.90" />
                    <SPLIT distance="150" swimtime="00:02:06.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="410" status="EXH" swimtime="00:01:06.54" resultid="6696" heatid="10709" lane="4" entrytime="00:01:04.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="404" status="EXH" swimtime="00:04:57.68" resultid="6697" heatid="10722" lane="0" entrytime="00:04:49.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                    <SPLIT distance="100" swimtime="00:01:09.49" />
                    <SPLIT distance="150" swimtime="00:01:47.58" />
                    <SPLIT distance="200" swimtime="00:02:25.48" />
                    <SPLIT distance="250" swimtime="00:03:03.87" />
                    <SPLIT distance="300" swimtime="00:03:41.97" />
                    <SPLIT distance="350" swimtime="00:04:20.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernanda" lastname="Vieira Gama" birthdate="2011-03-25" gender="F" nation="BRA" license="367948" swrid="5627396" athleteid="6698" externalid="367948">
              <RESULTS>
                <RESULT eventid="1147" points="357" status="EXH" swimtime="00:01:12.86" resultid="6699" heatid="10525" lane="8" />
                <RESULT eventid="1131" points="365" status="EXH" swimtime="00:06:09.91" resultid="6700" heatid="10519" lane="5" entrytime="00:06:08.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                    <SPLIT distance="100" swimtime="00:01:23.17" />
                    <SPLIT distance="150" swimtime="00:02:11.14" />
                    <SPLIT distance="200" swimtime="00:02:57.23" />
                    <SPLIT distance="250" swimtime="00:03:51.63" />
                    <SPLIT distance="300" swimtime="00:04:44.34" />
                    <SPLIT distance="350" swimtime="00:05:27.77" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 9:48)" eventid="1227" status="DSQ" swimtime="00:00:32.31" resultid="6701" heatid="10600" lane="2" />
                <RESULT eventid="1265" points="374" status="EXH" swimtime="00:02:55.02" resultid="6702" heatid="10642" lane="6" entrytime="00:02:50.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                    <SPLIT distance="100" swimtime="00:01:22.42" />
                    <SPLIT distance="150" swimtime="00:02:14.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="344" status="EXH" swimtime="00:05:35.85" resultid="6703" heatid="10714" lane="9" entrytime="00:05:29.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                    <SPLIT distance="100" swimtime="00:01:19.82" />
                    <SPLIT distance="150" swimtime="00:02:01.85" />
                    <SPLIT distance="200" swimtime="00:02:43.42" />
                    <SPLIT distance="250" swimtime="00:03:24.32" />
                    <SPLIT distance="300" swimtime="00:04:09.35" />
                    <SPLIT distance="350" swimtime="00:04:52.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="307" status="EXH" swimtime="00:01:21.76" resultid="6704" heatid="10701" lane="1" entrytime="00:01:20.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emanuel" lastname="Da Silva Scarantti" birthdate="2011-04-26" gender="M" nation="BRA" license="377367" athleteid="6733" externalid="377367">
              <RESULTS>
                <RESULT eventid="1123" points="307" status="EXH" swimtime="00:11:09.71" resultid="6734" heatid="10516" lane="7" entrytime="00:11:03.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.38" />
                    <SPLIT distance="100" swimtime="00:01:17.06" />
                    <SPLIT distance="150" swimtime="00:01:58.56" />
                    <SPLIT distance="200" swimtime="00:02:41.67" />
                    <SPLIT distance="250" swimtime="00:03:24.10" />
                    <SPLIT distance="300" swimtime="00:04:07.31" />
                    <SPLIT distance="350" swimtime="00:04:49.24" />
                    <SPLIT distance="400" swimtime="00:05:31.75" />
                    <SPLIT distance="450" swimtime="00:06:13.88" />
                    <SPLIT distance="500" swimtime="00:06:57.35" />
                    <SPLIT distance="550" swimtime="00:07:39.94" />
                    <SPLIT distance="600" swimtime="00:08:22.71" />
                    <SPLIT distance="650" swimtime="00:09:05.12" />
                    <SPLIT distance="700" swimtime="00:09:47.86" />
                    <SPLIT distance="750" swimtime="00:10:29.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="269" status="EXH" swimtime="00:03:14.17" resultid="6735" heatid="10489" lane="8" entrytime="00:03:10.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.01" />
                    <SPLIT distance="100" swimtime="00:01:32.28" />
                    <SPLIT distance="150" swimtime="00:02:24.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="264" swimtime="00:01:28.65" resultid="6736" heatid="10594" lane="0" entrytime="00:01:28.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="313" status="EXH" swimtime="00:02:30.10" resultid="6737" heatid="10667" lane="8" entrytime="00:02:30.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                    <SPLIT distance="100" swimtime="00:01:12.90" />
                    <SPLIT distance="150" swimtime="00:01:51.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="320" status="EXH" swimtime="00:05:21.52" resultid="6738" heatid="10719" lane="6" entrytime="00:05:25.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.13" />
                    <SPLIT distance="100" swimtime="00:01:14.41" />
                    <SPLIT distance="150" swimtime="00:01:54.96" />
                    <SPLIT distance="200" swimtime="00:02:36.17" />
                    <SPLIT distance="250" swimtime="00:03:17.53" />
                    <SPLIT distance="300" swimtime="00:03:59.78" />
                    <SPLIT distance="350" swimtime="00:04:41.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="253" status="EXH" swimtime="00:01:21.56" resultid="6739" heatid="10736" lane="1" entrytime="00:01:22.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Augusto Reitz" birthdate="2011-07-18" gender="M" nation="BRA" license="394878" athleteid="6775" externalid="394878">
              <RESULTS>
                <RESULT eventid="1087" points="221" status="EXH" swimtime="00:03:27.26" resultid="6776" heatid="10488" lane="1" entrytime="00:03:35.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.41" />
                    <SPLIT distance="100" swimtime="00:01:39.80" />
                    <SPLIT distance="150" swimtime="00:02:34.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="225" status="EXH" swimtime="00:01:16.26" resultid="6777" heatid="10537" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="209" status="EXH" swimtime="00:00:35.19" resultid="6778" heatid="10610" lane="2" />
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 9:28), Na volta dos 50m." eventid="1219" status="DSQ" swimtime="00:01:35.16" resultid="6779" heatid="10593" lane="0" entrytime="00:01:35.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="188" status="EXH" swimtime="00:03:18.90" resultid="6780" heatid="10646" lane="7" entrytime="00:03:16.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.78" />
                    <SPLIT distance="100" swimtime="00:01:43.21" />
                    <SPLIT distance="150" swimtime="00:02:36.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="251" status="EXH" swimtime="00:02:41.68" resultid="6781" heatid="10665" lane="4" entrytime="00:02:42.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                    <SPLIT distance="100" swimtime="00:01:18.15" />
                    <SPLIT distance="150" swimtime="00:02:00.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Menel Stahelin" birthdate="2006-01-25" gender="M" nation="BRA" license="298658" athleteid="6590" externalid="298658">
              <RESULTS>
                <RESULT eventid="1219" points="674" status="EXH" swimtime="00:01:04.85" resultid="6591" heatid="10599" lane="4" entrytime="00:01:03.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="532" status="EXH" swimtime="00:02:05.85" resultid="6592" heatid="10663" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.38" />
                    <SPLIT distance="100" swimtime="00:01:00.25" />
                    <SPLIT distance="150" swimtime="00:01:33.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Zayra" lastname="Thalya Maba" birthdate="2009-04-17" gender="F" nation="BRA" license="356024" swrid="5634815" athleteid="6649" externalid="356024">
              <RESULTS>
                <RESULT eventid="1079" points="327" status="EXH" swimtime="00:03:19.58" resultid="6650" heatid="10483" lane="9" entrytime="00:03:18.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.93" />
                    <SPLIT distance="100" swimtime="00:01:35.16" />
                    <SPLIT distance="150" swimtime="00:02:28.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="369" status="EXH" swimtime="00:06:08.51" resultid="6651" heatid="10519" lane="1" entrytime="00:06:17.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.82" />
                    <SPLIT distance="100" swimtime="00:01:20.84" />
                    <SPLIT distance="150" swimtime="00:02:09.53" />
                    <SPLIT distance="200" swimtime="00:02:57.33" />
                    <SPLIT distance="250" swimtime="00:03:48.08" />
                    <SPLIT distance="300" swimtime="00:04:40.13" />
                    <SPLIT distance="350" swimtime="00:05:26.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="333" status="EXH" swimtime="00:01:32.47" resultid="6652" heatid="10586" lane="0" entrytime="00:01:30.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="415" status="EXH" swimtime="00:02:49.02" resultid="6653" heatid="10642" lane="5" entrytime="00:02:49.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                    <SPLIT distance="100" swimtime="00:01:19.66" />
                    <SPLIT distance="150" swimtime="00:02:09.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="348" status="EXH" swimtime="00:02:39.42" resultid="6654" heatid="10653" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                    <SPLIT distance="100" swimtime="00:01:18.32" />
                    <SPLIT distance="150" swimtime="00:01:59.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="345" status="EXH" swimtime="00:01:18.65" resultid="6655" heatid="10701" lane="2" entrytime="00:01:18.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcus" lastname="Taylor Laraz" birthdate="2011-12-30" gender="M" nation="BRA" license="393411" athleteid="6761" externalid="393411">
              <RESULTS>
                <RESULT eventid="1087" points="199" status="EXH" swimtime="00:03:34.66" resultid="6762" heatid="10488" lane="7" entrytime="00:03:33.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.76" />
                    <SPLIT distance="100" swimtime="00:01:41.69" />
                    <SPLIT distance="150" swimtime="00:02:39.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="218" status="EXH" swimtime="00:01:17.09" resultid="6763" heatid="10539" lane="1" entrytime="00:01:15.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="194" status="EXH" swimtime="00:01:38.21" resultid="6764" heatid="10591" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="210" status="EXH" swimtime="00:03:11.65" resultid="6765" heatid="10646" lane="5" entrytime="00:03:11.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.07" />
                    <SPLIT distance="150" swimtime="00:02:28.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="231" status="EXH" swimtime="00:02:46.20" resultid="6766" heatid="10665" lane="1" entrytime="00:02:47.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="100" swimtime="00:01:19.52" />
                    <SPLIT distance="150" swimtime="00:02:04.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="195" status="EXH" swimtime="00:01:28.92" resultid="6767" heatid="10735" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Alves Dalzoto" birthdate="2012-09-14" gender="M" nation="BRA" license="381818" swrid="5748638" athleteid="6740" externalid="381818">
              <RESULTS>
                <RESULT eventid="1071" points="351" status="EXH" swimtime="00:02:38.55" resultid="6741" heatid="10477" lane="2" entrytime="00:02:38.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                    <SPLIT distance="100" swimtime="00:01:14.62" />
                    <SPLIT distance="150" swimtime="00:01:56.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="331" status="EXH" swimtime="00:01:07.05" resultid="6742" heatid="10543" lane="7" entrytime="00:01:07.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" status="WDR" swimtime="00:00:00.00" resultid="6743" heatid="10620" lane="8" entrytime="00:00:29.61" entrycourse="LCM" />
                <RESULT eventid="1273" status="WDR" swimtime="00:00:00.00" resultid="6744" heatid="10648" lane="9" entrytime="00:02:54.78" entrycourse="LCM" />
                <RESULT eventid="1341" status="WDR" swimtime="00:00:00.00" resultid="6745" heatid="10703" lane="2" />
                <RESULT eventid="1373" status="WDR" swimtime="00:00:00.00" resultid="6746" heatid="10738" lane="4" entrytime="00:01:13.61" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Hermenegildo" birthdate="2012-10-11" gender="F" nation="BRA" license="369477" swrid="5748687" athleteid="6726" externalid="369477">
              <RESULTS>
                <RESULT eventid="1079" points="391" status="EXH" swimtime="00:03:07.95" resultid="6727" heatid="10484" lane="8" entrytime="00:03:07.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.99" />
                    <SPLIT distance="100" swimtime="00:01:29.89" />
                    <SPLIT distance="150" swimtime="00:02:18.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="479" status="EXH" swimtime="00:02:37.30" resultid="6728" heatid="10473" lane="0" entrytime="00:02:39.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                    <SPLIT distance="100" swimtime="00:01:14.99" />
                    <SPLIT distance="150" swimtime="00:01:55.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="434" status="EXH" swimtime="00:05:49.06" resultid="6729" heatid="10520" lane="7" entrytime="00:05:50.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                    <SPLIT distance="100" swimtime="00:01:17.41" />
                    <SPLIT distance="150" swimtime="00:02:01.73" />
                    <SPLIT distance="200" swimtime="00:02:45.91" />
                    <SPLIT distance="250" swimtime="00:03:35.55" />
                    <SPLIT distance="300" swimtime="00:04:26.42" />
                    <SPLIT distance="350" swimtime="00:05:08.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="490" status="EXH" swimtime="00:02:39.91" resultid="6730" heatid="10644" lane="8" entrytime="00:02:41.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                    <SPLIT distance="100" swimtime="00:01:14.47" />
                    <SPLIT distance="150" swimtime="00:02:01.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="361" status="EXH" swimtime="00:01:17.49" resultid="6731" heatid="10699" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="464" status="EXH" swimtime="00:01:13.77" resultid="6732" heatid="10732" lane="8" entrytime="00:01:13.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Hillan Lisboa" birthdate="2007-05-08" gender="M" nation="BRA" license="327544" swrid="5634668" athleteid="6614" externalid="327544">
              <RESULTS>
                <RESULT eventid="1123" points="562" status="EXH" swimtime="00:09:07.83" resultid="6615" heatid="10513" lane="3" entrytime="00:08:56.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.08" />
                    <SPLIT distance="100" swimtime="00:01:05.03" />
                    <SPLIT distance="150" swimtime="00:01:38.74" />
                    <SPLIT distance="200" swimtime="00:02:12.77" />
                    <SPLIT distance="250" swimtime="00:02:47.63" />
                    <SPLIT distance="300" swimtime="00:03:22.04" />
                    <SPLIT distance="350" swimtime="00:03:56.52" />
                    <SPLIT distance="400" swimtime="00:04:31.14" />
                    <SPLIT distance="450" swimtime="00:05:06.33" />
                    <SPLIT distance="500" swimtime="00:05:41.29" />
                    <SPLIT distance="550" swimtime="00:06:16.58" />
                    <SPLIT distance="600" swimtime="00:06:51.55" />
                    <SPLIT distance="650" swimtime="00:07:26.80" />
                    <SPLIT distance="700" swimtime="00:08:01.40" />
                    <SPLIT distance="750" swimtime="00:08:35.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="480" status="EXH" swimtime="00:02:40.16" resultid="6616" heatid="10492" lane="8" entrytime="00:02:39.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.86" />
                    <SPLIT distance="100" swimtime="00:01:16.16" />
                    <SPLIT distance="150" swimtime="00:01:58.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="483" status="EXH" swimtime="00:05:08.92" resultid="6617" heatid="10523" lane="2" entrytime="00:05:00.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                    <SPLIT distance="100" swimtime="00:01:09.69" />
                    <SPLIT distance="150" swimtime="00:01:51.91" />
                    <SPLIT distance="200" swimtime="00:02:33.28" />
                    <SPLIT distance="250" swimtime="00:03:16.98" />
                    <SPLIT distance="300" swimtime="00:04:00.46" />
                    <SPLIT distance="350" swimtime="00:04:35.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="556" status="EXH" swimtime="00:17:38.38" resultid="6618" heatid="10635" lane="5" entrytime="00:17:15.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                    <SPLIT distance="100" swimtime="00:01:06.59" />
                    <SPLIT distance="150" swimtime="00:01:40.71" />
                    <SPLIT distance="200" swimtime="00:02:15.30" />
                    <SPLIT distance="250" swimtime="00:02:49.56" />
                    <SPLIT distance="300" swimtime="00:03:24.05" />
                    <SPLIT distance="350" swimtime="00:03:59.05" />
                    <SPLIT distance="400" swimtime="00:04:34.07" />
                    <SPLIT distance="450" swimtime="00:05:09.02" />
                    <SPLIT distance="500" swimtime="00:05:43.95" />
                    <SPLIT distance="550" swimtime="00:06:19.08" />
                    <SPLIT distance="600" swimtime="00:06:54.38" />
                    <SPLIT distance="650" swimtime="00:07:29.73" />
                    <SPLIT distance="700" swimtime="00:08:05.24" />
                    <SPLIT distance="750" swimtime="00:08:40.68" />
                    <SPLIT distance="800" swimtime="00:09:16.21" />
                    <SPLIT distance="850" swimtime="00:09:51.63" />
                    <SPLIT distance="900" swimtime="00:10:27.52" />
                    <SPLIT distance="950" swimtime="00:11:03.77" />
                    <SPLIT distance="1000" swimtime="00:11:39.96" />
                    <SPLIT distance="1050" swimtime="00:12:16.06" />
                    <SPLIT distance="1100" swimtime="00:12:52.43" />
                    <SPLIT distance="1150" swimtime="00:13:28.89" />
                    <SPLIT distance="1200" swimtime="00:14:05.09" />
                    <SPLIT distance="1250" swimtime="00:14:41.18" />
                    <SPLIT distance="1300" swimtime="00:15:17.41" />
                    <SPLIT distance="1350" swimtime="00:15:53.30" />
                    <SPLIT distance="1400" swimtime="00:16:28.55" />
                    <SPLIT distance="1450" swimtime="00:17:03.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="442" status="EXH" swimtime="00:02:29.59" resultid="6619" heatid="10652" lane="2" entrytime="00:02:19.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                    <SPLIT distance="100" swimtime="00:01:12.64" />
                    <SPLIT distance="150" swimtime="00:01:54.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="561" status="EXH" swimtime="00:04:26.74" resultid="6620" heatid="10724" lane="6" entrytime="00:04:19.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.13" />
                    <SPLIT distance="100" swimtime="00:01:02.26" />
                    <SPLIT distance="150" swimtime="00:01:35.41" />
                    <SPLIT distance="200" swimtime="00:02:09.34" />
                    <SPLIT distance="250" swimtime="00:02:43.01" />
                    <SPLIT distance="300" swimtime="00:03:17.78" />
                    <SPLIT distance="350" swimtime="00:03:52.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Menine Schneider" birthdate="2012-12-05" gender="M" nation="BRA" license="393406" athleteid="6754" externalid="393406">
              <RESULTS>
                <RESULT eventid="1087" points="194" status="EXH" swimtime="00:03:36.57" resultid="6755" heatid="10488" lane="8" entrytime="00:03:41.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.67" />
                    <SPLIT distance="100" swimtime="00:01:43.00" />
                    <SPLIT distance="150" swimtime="00:02:40.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="235" status="EXH" swimtime="00:00:42.00" resultid="6756" heatid="10571" lane="2" entrytime="00:00:42.89" entrycourse="LCM" />
                <RESULT eventid="1155" points="248" status="EXH" swimtime="00:01:13.84" resultid="6757" heatid="10540" lane="9" entrytime="00:01:14.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="193" status="EXH" swimtime="00:01:38.38" resultid="6758" heatid="10592" lane="5" entrytime="00:01:38.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.21" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 8.3 - Movimento alternado das pernas ou pés.  (Horário: 16:32), Na volta dos 50m (Borboleta, Medley Individual)." eventid="1273" status="DSQ" swimtime="00:03:30.15" resultid="6759" heatid="10646" lane="8" entrytime="00:03:25.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:52.28" />
                    <SPLIT distance="150" swimtime="00:02:48.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="228" status="EXH" swimtime="00:02:46.93" resultid="6760" heatid="10665" lane="7" entrytime="00:02:45.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                    <SPLIT distance="100" swimtime="00:01:21.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Matejczyk" birthdate="2011-07-04" gender="M" nation="BRA" license="399784" athleteid="6789" externalid="399784">
              <RESULTS>
                <RESULT eventid="1071" points="367" status="EXH" swimtime="00:02:36.24" resultid="6790" heatid="10477" lane="3" entrytime="00:02:36.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                    <SPLIT distance="100" swimtime="00:01:13.31" />
                    <SPLIT distance="150" swimtime="00:01:54.78" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 18:10)" eventid="1155" status="DSQ" swimtime="00:01:02.61" resultid="6791" heatid="10545" lane="3" entrytime="00:01:04.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="394" status="EXH" swimtime="00:00:28.50" resultid="6792" heatid="10621" lane="2" entrytime="00:00:28.61" entrycourse="LCM" />
                <RESULT eventid="1219" points="296" status="EXH" swimtime="00:01:25.28" resultid="6793" heatid="10594" lane="9" entrytime="00:01:29.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="396" status="EXH" swimtime="00:02:18.86" resultid="6794" heatid="10669" lane="7" entrytime="00:02:19.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                    <SPLIT distance="100" swimtime="00:01:05.44" />
                    <SPLIT distance="150" swimtime="00:01:42.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="395" status="EXH" swimtime="00:04:59.73" resultid="6795" heatid="10718" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                    <SPLIT distance="100" swimtime="00:01:11.18" />
                    <SPLIT distance="150" swimtime="00:01:50.54" />
                    <SPLIT distance="200" swimtime="00:02:29.09" />
                    <SPLIT distance="250" swimtime="00:03:07.59" />
                    <SPLIT distance="300" swimtime="00:03:46.35" />
                    <SPLIT distance="350" swimtime="00:04:24.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joanna" lastname="Beatriz Rossi" birthdate="2006-03-01" gender="F" nation="BRA" license="318797" athleteid="6593" externalid="318797">
              <RESULTS>
                <RESULT eventid="1079" points="552" status="EXH" swimtime="00:02:47.61" resultid="6594" heatid="10486" lane="5" entrytime="00:02:45.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.65" />
                    <SPLIT distance="100" swimtime="00:01:19.09" />
                    <SPLIT distance="150" swimtime="00:02:03.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="538" status="EXH" swimtime="00:00:35.85" resultid="6595" heatid="10565" lane="5" entrytime="00:00:35.29" entrycourse="LCM" />
                <RESULT eventid="1147" points="653" status="EXH" swimtime="00:00:59.58" resultid="6596" heatid="10534" lane="5" entrytime="00:01:00.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="573" status="EXH" swimtime="00:01:17.19" resultid="6597" heatid="10589" lane="5" entrytime="00:01:14.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="627" status="EXH" swimtime="00:02:27.30" resultid="6598" heatid="10644" lane="4" entrytime="00:02:25.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.47" />
                    <SPLIT distance="100" swimtime="00:01:09.58" />
                    <SPLIT distance="150" swimtime="00:01:52.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="587" status="EXH" swimtime="00:01:05.90" resultid="6599" heatid="10699" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Gabriel Do Prado" birthdate="2010-01-05" gender="M" nation="BRA" license="367935" swrid="5588710" athleteid="6677" externalid="367935">
              <RESULTS>
                <RESULT eventid="1071" points="442" status="EXH" swimtime="00:02:26.88" resultid="6678" heatid="10479" lane="0" entrytime="00:02:26.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                    <SPLIT distance="100" swimtime="00:01:11.12" />
                    <SPLIT distance="150" swimtime="00:01:48.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="559" status="EXH" swimtime="00:00:56.31" resultid="6679" heatid="10551" lane="2" entrytime="00:00:55.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="487" status="EXH" swimtime="00:02:24.85" resultid="6680" heatid="10651" lane="4" entrytime="00:02:22.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.92" />
                    <SPLIT distance="100" swimtime="00:01:05.89" />
                    <SPLIT distance="150" swimtime="00:01:49.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="511" status="EXH" swimtime="00:02:07.52" resultid="6681" heatid="10672" lane="4" entrytime="00:02:08.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.36" />
                    <SPLIT distance="100" swimtime="00:01:01.24" />
                    <SPLIT distance="150" swimtime="00:01:34.11" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 9:25), Na volta dos 50m." eventid="1341" status="DSQ" swimtime="00:01:05.41" resultid="6682" heatid="10710" lane="0" entrytime="00:01:04.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="475" status="EXH" swimtime="00:01:06.13" resultid="6683" heatid="10742" lane="9" entrytime="00:01:04.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Lennert" birthdate="2007-10-04" gender="M" nation="BRA" license="327536" swrid="5634686" athleteid="6600" externalid="327536">
              <RESULTS>
                <RESULT eventid="1103" points="626" status="EXH" swimtime="00:00:26.03" resultid="6601" heatid="10508" lane="3" entrytime="00:00:26.30" entrycourse="LCM" />
                <RESULT eventid="1155" points="615" status="EXH" swimtime="00:00:54.55" resultid="6602" heatid="10552" lane="9" entrytime="00:00:54.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="593" status="EXH" swimtime="00:00:24.88" resultid="6603" heatid="10627" lane="3" entrytime="00:00:25.18" entrycourse="LCM" />
                <RESULT eventid="1273" points="562" status="EXH" swimtime="00:02:18.12" resultid="6604" heatid="10652" lane="6" entrytime="00:02:18.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                    <SPLIT distance="100" swimtime="00:01:04.26" />
                    <SPLIT distance="150" swimtime="00:01:47.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="620" status="EXH" swimtime="00:00:57.98" resultid="6605" heatid="10711" lane="3" entrytime="00:00:58.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="557" status="EXH" swimtime="00:01:02.71" resultid="6606" heatid="10734" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Gonçalves Sguário" birthdate="2009-04-27" gender="M" nation="BRA" license="369471" swrid="5634654" athleteid="6719" externalid="369471">
              <RESULTS>
                <RESULT eventid="1071" points="449" status="EXH" swimtime="00:02:26.13" resultid="6720" heatid="10480" lane="9" entrytime="00:02:24.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                    <SPLIT distance="100" swimtime="00:01:10.24" />
                    <SPLIT distance="150" swimtime="00:01:48.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="563" status="EXH" swimtime="00:00:56.18" resultid="6721" heatid="10551" lane="3" entrytime="00:00:55.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="548" status="EXH" swimtime="00:00:25.55" resultid="6722" heatid="10626" lane="2" entrytime="00:00:25.82" entrycourse="LCM" />
                <RESULT eventid="1273" points="434" status="EXH" swimtime="00:02:30.57" resultid="6723" heatid="10650" lane="3" entrytime="00:02:31.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                    <SPLIT distance="100" swimtime="00:01:11.07" />
                    <SPLIT distance="150" swimtime="00:01:57.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="482" status="EXH" swimtime="00:02:10.07" resultid="6724" heatid="10673" lane="9" entrytime="00:02:07.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                    <SPLIT distance="100" swimtime="00:01:02.18" />
                    <SPLIT distance="150" swimtime="00:01:36.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="524" status="EXH" swimtime="00:01:03.97" resultid="6725" heatid="10741" lane="3" entrytime="00:01:04.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Vitor Ivaldo Da Costa Pereira" birthdate="2010-07-06" gender="M" nation="BRA" license="356025" swrid="5588956" athleteid="6656" externalid="356025">
              <RESULTS>
                <RESULT eventid="1087" points="547" status="EXH" swimtime="00:02:33.41" resultid="6657" heatid="10492" lane="6" entrytime="00:02:31.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                    <SPLIT distance="100" swimtime="00:01:13.93" />
                    <SPLIT distance="150" swimtime="00:01:54.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="471" status="EXH" swimtime="00:05:11.51" resultid="6658" heatid="10523" lane="7" entrytime="00:05:04.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.85" />
                    <SPLIT distance="100" swimtime="00:01:10.41" />
                    <SPLIT distance="150" swimtime="00:01:52.80" />
                    <SPLIT distance="200" swimtime="00:02:34.82" />
                    <SPLIT distance="250" swimtime="00:03:16.77" />
                    <SPLIT distance="300" swimtime="00:03:58.63" />
                    <SPLIT distance="350" swimtime="00:04:35.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="492" status="EXH" swimtime="00:01:12.05" resultid="6659" heatid="10598" lane="3" entrytime="00:01:10.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="479" status="EXH" swimtime="00:02:25.70" resultid="6660" heatid="10652" lane="0" entrytime="00:02:22.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                    <SPLIT distance="100" swimtime="00:01:12.61" />
                    <SPLIT distance="150" swimtime="00:01:52.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="408" status="EXH" swimtime="00:01:06.64" resultid="6661" heatid="10709" lane="1" entrytime="00:01:06.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="406" status="EXH" swimtime="00:01:09.63" resultid="6662" heatid="10734" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Paulus Negherbon" birthdate="2009-10-01" gender="F" nation="BRA" license="347400" swrid="5634752" athleteid="6635" externalid="347400">
              <RESULTS>
                <RESULT eventid="1063" points="532" status="EXH" swimtime="00:02:31.92" resultid="6636" heatid="10473" lane="5" entrytime="00:02:31.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.97" />
                    <SPLIT distance="100" swimtime="00:01:12.66" />
                    <SPLIT distance="150" swimtime="00:01:52.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="493" status="EXH" swimtime="00:02:34.09" resultid="6637" heatid="10554" lane="5" entrytime="00:02:30.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.17" />
                    <SPLIT distance="100" swimtime="00:01:11.28" />
                    <SPLIT distance="150" swimtime="00:01:52.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="523" status="EXH" swimtime="00:05:28.09" resultid="6638" heatid="10520" lane="4" entrytime="00:05:21.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                    <SPLIT distance="100" swimtime="00:01:10.49" />
                    <SPLIT distance="150" swimtime="00:01:51.56" />
                    <SPLIT distance="200" swimtime="00:02:32.41" />
                    <SPLIT distance="250" swimtime="00:03:21.40" />
                    <SPLIT distance="300" swimtime="00:04:10.47" />
                    <SPLIT distance="350" swimtime="00:04:49.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="527" status="EXH" swimtime="00:02:36.08" resultid="6639" heatid="10644" lane="5" entrytime="00:02:33.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                    <SPLIT distance="100" swimtime="00:01:11.67" />
                    <SPLIT distance="150" swimtime="00:01:59.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="477" status="EXH" swimtime="00:02:23.62" resultid="6640" heatid="10660" lane="7" entrytime="00:02:18.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                    <SPLIT distance="100" swimtime="00:01:09.27" />
                    <SPLIT distance="150" swimtime="00:01:46.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="531" status="EXH" swimtime="00:01:10.53" resultid="6641" heatid="10726" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Zimmermann Da Silva" birthdate="2010-05-10" gender="F" nation="BRA" license="362474" swrid="5588673" athleteid="6670" externalid="362474">
              <RESULTS>
                <RESULT eventid="1079" points="479" status="EXH" swimtime="00:02:55.73" resultid="6671" heatid="10485" lane="3" entrytime="00:02:57.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.06" />
                    <SPLIT distance="100" swimtime="00:01:24.84" />
                    <SPLIT distance="150" swimtime="00:02:11.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="388" status="EXH" swimtime="00:02:46.96" resultid="6672" heatid="10554" lane="3" entrytime="00:02:42.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.45" />
                    <SPLIT distance="100" swimtime="00:01:19.25" />
                    <SPLIT distance="150" swimtime="00:02:04.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="439" status="EXH" swimtime="00:01:24.38" resultid="6673" heatid="10588" lane="3" entrytime="00:01:21.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="442" status="EXH" swimtime="00:02:45.55" resultid="6674" heatid="10644" lane="7" entrytime="00:02:40.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.21" />
                    <SPLIT distance="100" swimtime="00:01:20.20" />
                    <SPLIT distance="150" swimtime="00:02:08.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="449" status="EXH" swimtime="00:02:26.50" resultid="6675" heatid="10660" lane="9" entrytime="00:02:20.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="100" swimtime="00:01:11.76" />
                    <SPLIT distance="150" swimtime="00:01:49.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="480" status="EXH" swimtime="00:05:00.54" resultid="6676" heatid="10716" lane="6" entrytime="00:04:57.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                    <SPLIT distance="100" swimtime="00:01:12.55" />
                    <SPLIT distance="150" swimtime="00:01:50.52" />
                    <SPLIT distance="200" swimtime="00:02:28.91" />
                    <SPLIT distance="250" swimtime="00:03:06.44" />
                    <SPLIT distance="300" swimtime="00:03:44.44" />
                    <SPLIT distance="350" swimtime="00:04:23.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Kayan Fontineli" birthdate="2011-09-05" gender="M" nation="BRA" license="393415" athleteid="6768" externalid="393415">
              <RESULTS>
                <RESULT eventid="1155" points="430" status="EXH" swimtime="00:01:01.44" resultid="6769" heatid="10547" lane="2" entrytime="00:01:01.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="426" status="EXH" swimtime="00:00:27.77" resultid="6770" heatid="10623" lane="8" entrytime="00:00:27.77" entrycourse="LCM" />
                <RESULT eventid="1273" points="361" status="EXH" swimtime="00:02:40.09" resultid="6771" heatid="10649" lane="1" entrytime="00:02:43.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                    <SPLIT distance="100" swimtime="00:01:17.21" />
                    <SPLIT distance="150" swimtime="00:02:03.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="412" status="EXH" swimtime="00:02:16.99" resultid="6772" heatid="10670" lane="4" entrytime="00:02:16.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                    <SPLIT distance="100" swimtime="00:01:06.02" />
                    <SPLIT distance="150" swimtime="00:01:41.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="388" status="EXH" swimtime="00:05:01.49" resultid="6773" heatid="10721" lane="7" entrytime="00:04:55.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                    <SPLIT distance="100" swimtime="00:01:09.89" />
                    <SPLIT distance="150" swimtime="00:01:48.34" />
                    <SPLIT distance="200" swimtime="00:02:26.96" />
                    <SPLIT distance="250" swimtime="00:03:05.46" />
                    <SPLIT distance="300" swimtime="00:03:44.00" />
                    <SPLIT distance="350" swimtime="00:04:22.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="274" status="EXH" swimtime="00:01:19.40" resultid="6774" heatid="10737" lane="7" entrytime="00:01:18.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Richard" lastname="Fiorelli" birthdate="2011-01-26" gender="M" nation="BRA" license="385730" swrid="5684554" athleteid="6747" externalid="385730">
              <RESULTS>
                <RESULT eventid="1071" points="326" status="EXH" swimtime="00:02:42.48" resultid="6748" heatid="10477" lane="7" entrytime="00:02:41.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                    <SPLIT distance="100" swimtime="00:01:16.57" />
                    <SPLIT distance="150" swimtime="00:01:59.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="374" status="EXH" swimtime="00:01:04.38" resultid="6749" heatid="10545" lane="8" entrytime="00:01:04.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="370" status="EXH" swimtime="00:00:29.12" resultid="6750" heatid="10621" lane="9" entrytime="00:00:29.01" entrycourse="LCM" />
                <RESULT eventid="1273" points="311" status="EXH" swimtime="00:02:48.11" resultid="6751" heatid="10648" lane="6" entrytime="00:02:50.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                    <SPLIT distance="100" swimtime="00:01:16.53" />
                    <SPLIT distance="150" swimtime="00:02:08.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="309" status="EXH" swimtime="00:02:30.74" resultid="6752" heatid="10668" lane="9" entrytime="00:02:26.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                    <SPLIT distance="100" swimtime="00:01:09.02" />
                    <SPLIT distance="150" swimtime="00:01:49.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="351" status="EXH" swimtime="00:01:13.09" resultid="6753" heatid="10738" lane="6" entrytime="00:01:14.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Celestino Da Silva" birthdate="2007-01-17" gender="M" nation="BRA" license="327540" swrid="5634558" athleteid="6607" externalid="327540">
              <RESULTS>
                <RESULT eventid="1103" points="481" status="EXH" swimtime="00:00:28.42" resultid="6608" heatid="10507" lane="6" entrytime="00:00:28.30" entrycourse="LCM" />
                <RESULT eventid="1187" points="474" status="EXH" swimtime="00:00:33.27" resultid="6609" heatid="10574" lane="5" entrytime="00:00:32.47" entrycourse="LCM" />
                <RESULT eventid="1155" points="509" status="EXH" swimtime="00:00:58.11" resultid="6610" heatid="10549" lane="8" entrytime="00:00:59.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="439" status="EXH" swimtime="00:01:14.80" resultid="6611" heatid="10597" lane="4" entrytime="00:01:13.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 6.4 - A virada não foi iniciada após a conclusão do movimento de braço, após sair da posição de costas.  (Horário: 16:32), Na volta dos 100m (Costas, Medley Individual)." eventid="1273" status="DSQ" swimtime="00:02:29.46" resultid="6612" heatid="10646" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                    <SPLIT distance="100" swimtime="00:01:10.95" />
                    <SPLIT distance="150" swimtime="00:01:55.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="461" status="EXH" swimtime="00:01:03.99" resultid="6613" heatid="10710" lane="2" entrytime="00:01:02.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2539" nation="BRA" region="PR" clubid="7521" swrid="93771" name="Círculo Militar Do Paraná" shortname="Círculo Militar">
          <ATHLETES>
            <ATHLETE firstname="Vicente" lastname="Bileski" birthdate="2011-06-29" gender="M" nation="BRA" license="406950" swrid="5717248" athleteid="7546" externalid="406950">
              <RESULTS>
                <RESULT eventid="1103" points="293" swimtime="00:00:33.50" resultid="7547" heatid="10504" lane="1" entrytime="00:00:34.00" entrycourse="LCM" />
                <RESULT eventid="1155" points="330" swimtime="00:01:07.11" resultid="7548" heatid="10540" lane="2" entrytime="00:01:13.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="320" swimtime="00:00:30.56" resultid="7549" heatid="10617" lane="7" entrytime="00:00:31.16" entrycourse="LCM" />
                <RESULT eventid="1273" points="261" swimtime="00:02:58.23" resultid="7550" heatid="10646" lane="6" entrytime="00:03:11.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                    <SPLIT distance="100" swimtime="00:01:22.03" />
                    <SPLIT distance="150" swimtime="00:02:18.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Maria Romanelli" birthdate="2011-04-18" gender="F" nation="BRA" license="378335" swrid="5588803" athleteid="7535" externalid="378335">
              <RESULTS>
                <RESULT eventid="1095" points="239" swimtime="00:00:39.32" resultid="7536" heatid="10496" lane="2" entrytime="00:00:37.40" entrycourse="LCM" />
                <RESULT eventid="1227" points="384" swimtime="00:00:32.47" resultid="7537" heatid="10605" lane="0" entrytime="00:00:31.52" entrycourse="LCM" />
                <RESULT eventid="1297" points="314" swimtime="00:00:39.51" resultid="7538" heatid="10678" lane="4" entrytime="00:00:40.02" entrycourse="LCM" />
                <RESULT eventid="1265" points="278" swimtime="00:03:13.19" resultid="7539" heatid="10639" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                    <SPLIT distance="100" swimtime="00:01:32.37" />
                    <SPLIT distance="150" swimtime="00:02:34.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="281" swimtime="00:01:27.22" resultid="7540" heatid="10728" lane="5" entrytime="00:01:26.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernando" lastname="Jun Melo Ogima" birthdate="2006-07-05" gender="M" nation="BRA" license="378332" swrid="5622284" athleteid="7529" externalid="378332">
              <RESULTS>
                <RESULT eventid="1103" points="398" swimtime="00:00:30.26" resultid="7530" heatid="10506" lane="9" entrytime="00:00:30.96" entrycourse="LCM" />
                <RESULT eventid="1187" points="347" swimtime="00:00:36.92" resultid="7531" heatid="10568" lane="2" />
                <RESULT eventid="1219" points="293" swimtime="00:01:25.58" resultid="7532" heatid="10594" lane="2" entrytime="00:01:27.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="297" swimtime="00:02:50.84" resultid="7533" heatid="10648" lane="7" entrytime="00:02:51.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.99" />
                    <SPLIT distance="100" swimtime="00:01:18.22" />
                    <SPLIT distance="150" swimtime="00:02:08.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="239" swimtime="00:01:19.58" resultid="7534" heatid="10707" lane="9" entrytime="00:01:15.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Flavia" lastname="Scheffler Souza" birthdate="2010-09-14" gender="F" nation="BRA" license="417278" swrid="5757095" athleteid="7553" externalid="417278">
              <RESULTS>
                <RESULT eventid="1147" points="425" swimtime="00:01:08.73" resultid="7554" heatid="10530" lane="0" entrytime="00:01:08.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="381" swimtime="00:02:34.73" resultid="7555" heatid="10656" lane="2" entrytime="00:02:33.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                    <SPLIT distance="100" swimtime="00:01:11.44" />
                    <SPLIT distance="150" swimtime="00:01:52.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Manocchio" birthdate="2011-07-28" gender="M" nation="BRA" license="384916" swrid="5588573" athleteid="7541" externalid="384916">
              <RESULTS>
                <RESULT eventid="1155" points="390" swimtime="00:01:03.48" resultid="7542" heatid="10546" lane="8" entrytime="00:01:03.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="395" swimtime="00:00:28.48" resultid="7543" heatid="10621" lane="5" entrytime="00:00:28.43" entrycourse="LCM" />
                <RESULT eventid="1289" points="361" swimtime="00:02:23.18" resultid="7544" heatid="10669" lane="8" entrytime="00:02:20.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.79" />
                    <SPLIT distance="100" swimtime="00:01:07.29" />
                    <SPLIT distance="150" swimtime="00:01:45.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" status="DNS" swimtime="00:00:00.00" resultid="7545" heatid="10719" lane="5" entrytime="00:05:18.44" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Vieira De Macedo Brasil" birthdate="2009-12-19" gender="F" nation="BRA" license="344143" swrid="5622311" athleteid="7522" externalid="344143">
              <RESULTS>
                <RESULT eventid="1179" points="330" swimtime="00:00:42.17" resultid="7523" heatid="10563" lane="2" entrytime="00:00:41.42" entrycourse="LCM" />
                <RESULT eventid="1147" points="451" swimtime="00:01:07.38" resultid="7524" heatid="10530" lane="8" entrytime="00:01:08.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="406" swimtime="00:00:31.86" resultid="7525" heatid="10605" lane="2" entrytime="00:00:31.41" entrycourse="LCM" />
                <RESULT eventid="1211" points="306" swimtime="00:01:35.07" resultid="7526" heatid="10585" lane="3" entrytime="00:01:31.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="309" swimtime="00:03:06.51" resultid="7527" heatid="10640" lane="3" entrytime="00:03:12.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.37" />
                    <SPLIT distance="100" swimtime="00:01:35.44" />
                    <SPLIT distance="150" swimtime="00:02:28.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="363" swimtime="00:05:29.71" resultid="7528" heatid="10713" lane="3" entrytime="00:05:34.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                    <SPLIT distance="100" swimtime="00:01:19.79" />
                    <SPLIT distance="150" swimtime="00:02:03.88" />
                    <SPLIT distance="200" swimtime="00:02:48.72" />
                    <SPLIT distance="250" swimtime="00:03:29.83" />
                    <SPLIT distance="300" swimtime="00:04:11.05" />
                    <SPLIT distance="350" swimtime="00:04:51.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Oliveira Martini" birthdate="2008-10-31" gender="M" nation="BRA" license="406953" swrid="5717285" athleteid="7551" externalid="406953">
              <RESULTS>
                <RESULT eventid="1289" points="371" swimtime="00:02:21.84" resultid="7552" heatid="10668" lane="3" entrytime="00:02:21.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.20" />
                    <SPLIT distance="100" swimtime="00:01:07.69" />
                    <SPLIT distance="150" swimtime="00:01:45.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanna" lastname="Devitte Piegel" birthdate="2010-07-15" gender="F" nation="BRA" license="423469" athleteid="7556" externalid="423469">
              <RESULTS>
                <RESULT eventid="1227" points="112" swimtime="00:00:48.88" resultid="7557" heatid="10600" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16131" nation="BRA" region="PR" clubid="8503" swrid="93766" name="Associação Nadar Colombo" shortname="Equipe Nadar">
          <ATHLETES>
            <ATHLETE firstname="Nicole" lastname="Videira" birthdate="2010-08-10" gender="F" nation="BRA" license="421430" swrid="5811242" athleteid="8533" externalid="421430">
              <RESULTS>
                <RESULT eventid="1079" points="185" swimtime="00:04:01.04" resultid="8534" heatid="10482" lane="8" entrytime="00:04:03.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.15" />
                    <SPLIT distance="100" swimtime="00:01:53.68" />
                    <SPLIT distance="150" swimtime="00:02:58.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="223" swimtime="00:00:48.06" resultid="8535" heatid="10560" lane="4" />
                <RESULT eventid="1227" points="267" swimtime="00:00:36.64" resultid="8536" heatid="10602" lane="0" entrytime="00:00:36.93" entrycourse="LCM" />
                <RESULT eventid="1211" points="204" swimtime="00:01:48.79" resultid="8537" heatid="10583" lane="4" entrytime="00:01:51.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Santos Poli" birthdate="2010-02-19" gender="M" nation="BRA" license="414563" swrid="5755378" athleteid="8529" externalid="414563">
              <RESULTS>
                <RESULT eventid="1103" points="409" swimtime="00:00:30.00" resultid="8530" heatid="10506" lane="7" entrytime="00:00:30.48" entrycourse="LCM" />
                <RESULT eventid="1235" points="398" swimtime="00:00:28.41" resultid="8531" heatid="10618" lane="7" entrytime="00:00:30.68" entrycourse="LCM" />
                <RESULT eventid="1341" points="318" swimtime="00:01:12.40" resultid="8532" heatid="10707" lane="6" entrytime="00:01:12.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tayna" lastname="Macedo Gabardo" birthdate="2012-12-01" gender="F" nation="BRA" license="406704" swrid="5717281" athleteid="8523" externalid="406704">
              <RESULTS>
                <RESULT eventid="1063" points="239" swimtime="00:03:18.27" resultid="8524" heatid="10469" lane="4" entrytime="00:03:23.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="247" swimtime="00:01:22.41" resultid="8525" heatid="10527" lane="9" entrytime="00:01:18.58" entrycourse="LCM" />
                <RESULT eventid="1227" points="290" swimtime="00:00:35.65" resultid="8526" heatid="10602" lane="2" entrytime="00:00:35.53" entrycourse="LCM" />
                <RESULT eventid="1297" points="275" swimtime="00:00:41.29" resultid="8527" heatid="10678" lane="6" entrytime="00:00:40.94" entrycourse="LCM" />
                <RESULT eventid="1365" points="245" swimtime="00:01:31.19" resultid="8528" heatid="10727" lane="5" entrytime="00:01:30.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Glir" birthdate="2010-07-01" gender="M" nation="BRA" license="406701" swrid="5717266" athleteid="8518" externalid="406701">
              <RESULTS>
                <RESULT eventid="1187" points="235" swimtime="00:00:42.05" resultid="8519" heatid="10571" lane="3" entrytime="00:00:41.05" entrycourse="LCM" />
                <RESULT eventid="1155" points="407" swimtime="00:01:02.61" resultid="8520" heatid="10547" lane="9" entrytime="00:01:02.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="379" swimtime="00:00:28.89" resultid="8521" heatid="10622" lane="3" entrytime="00:00:27.98" entrycourse="LCM" />
                <RESULT eventid="1219" status="DNS" swimtime="00:00:00.00" resultid="8522" heatid="10593" lane="1" entrytime="00:01:32.65" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Rafael D Agostin Batistao" birthdate="2008-05-13" gender="M" nation="BRA" license="384738" swrid="5622300" athleteid="8504" externalid="384738">
              <RESULTS>
                <RESULT eventid="1187" points="341" swimtime="00:00:37.12" resultid="8505" heatid="10573" lane="1" entrytime="00:00:36.11" entrycourse="LCM" />
                <RESULT eventid="1235" points="362" swimtime="00:00:29.32" resultid="8506" heatid="10618" lane="1" entrytime="00:00:30.70" entrycourse="LCM" />
                <RESULT eventid="1219" points="342" swimtime="00:01:21.31" resultid="8507" heatid="10595" lane="6" entrytime="00:01:22.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lara" lastname="Carvalho Ezaki" birthdate="2011-10-20" gender="F" nation="BRA" license="399927" swrid="5652882" athleteid="8512" externalid="399927">
              <RESULTS>
                <RESULT eventid="1079" points="290" swimtime="00:03:27.68" resultid="8513" heatid="10482" lane="7" entrytime="00:03:30.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.65" />
                    <SPLIT distance="100" swimtime="00:01:42.40" />
                    <SPLIT distance="150" swimtime="00:02:37.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="169" swimtime="00:03:40.10" resultid="8514" heatid="10553" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.47" />
                    <SPLIT distance="100" swimtime="00:01:44.51" />
                    <SPLIT distance="150" swimtime="00:02:44.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="289" swimtime="00:01:36.90" resultid="8515" heatid="10584" lane="6" entrytime="00:01:37.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="306" swimtime="00:03:07.14" resultid="8516" heatid="10640" lane="2" entrytime="00:03:14.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.81" />
                    <SPLIT distance="150" swimtime="00:02:28.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="211" swimtime="00:01:32.66" resultid="8517" heatid="10699" lane="4" entrytime="00:01:45.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Luiz Sartori" birthdate="2008-04-07" gender="M" nation="BRA" license="384742" swrid="5622287" athleteid="8508" externalid="384742">
              <RESULTS>
                <RESULT eventid="1123" points="316" swimtime="00:11:03.21" resultid="8509" heatid="10517" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                    <SPLIT distance="100" swimtime="00:01:15.11" />
                    <SPLIT distance="150" swimtime="00:01:56.76" />
                    <SPLIT distance="200" swimtime="00:02:38.58" />
                    <SPLIT distance="250" swimtime="00:03:21.16" />
                    <SPLIT distance="300" swimtime="00:04:03.89" />
                    <SPLIT distance="350" swimtime="00:04:47.14" />
                    <SPLIT distance="400" swimtime="00:05:30.46" />
                    <SPLIT distance="450" swimtime="00:06:13.10" />
                    <SPLIT distance="500" swimtime="00:06:56.28" />
                    <SPLIT distance="550" swimtime="00:07:38.43" />
                    <SPLIT distance="600" swimtime="00:08:20.82" />
                    <SPLIT distance="650" swimtime="00:09:01.77" />
                    <SPLIT distance="700" swimtime="00:09:43.40" />
                    <SPLIT distance="750" swimtime="00:10:23.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="309" swimtime="00:21:27.19" resultid="8510" heatid="10637" lane="0" entrytime="00:21:44.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.69" />
                    <SPLIT distance="100" swimtime="00:01:17.92" />
                    <SPLIT distance="150" swimtime="00:02:00.38" />
                    <SPLIT distance="200" swimtime="00:02:43.59" />
                    <SPLIT distance="250" swimtime="00:03:27.04" />
                    <SPLIT distance="300" swimtime="00:04:10.84" />
                    <SPLIT distance="350" swimtime="00:04:54.76" />
                    <SPLIT distance="400" swimtime="00:05:38.39" />
                    <SPLIT distance="450" swimtime="00:06:22.23" />
                    <SPLIT distance="500" swimtime="00:07:05.06" />
                    <SPLIT distance="550" swimtime="00:07:48.29" />
                    <SPLIT distance="600" swimtime="00:08:32.10" />
                    <SPLIT distance="650" swimtime="00:09:15.73" />
                    <SPLIT distance="700" swimtime="00:09:59.59" />
                    <SPLIT distance="750" swimtime="00:10:43.45" />
                    <SPLIT distance="800" swimtime="00:11:27.09" />
                    <SPLIT distance="850" swimtime="00:12:10.55" />
                    <SPLIT distance="900" swimtime="00:12:54.34" />
                    <SPLIT distance="950" swimtime="00:13:37.89" />
                    <SPLIT distance="1000" swimtime="00:14:21.47" />
                    <SPLIT distance="1050" swimtime="00:15:04.04" />
                    <SPLIT distance="1100" swimtime="00:15:47.26" />
                    <SPLIT distance="1150" swimtime="00:16:30.18" />
                    <SPLIT distance="1200" swimtime="00:17:13.40" />
                    <SPLIT distance="1250" swimtime="00:17:56.46" />
                    <SPLIT distance="1300" swimtime="00:18:39.72" />
                    <SPLIT distance="1350" swimtime="00:19:22.22" />
                    <SPLIT distance="1400" swimtime="00:20:05.33" />
                    <SPLIT distance="1450" swimtime="00:20:47.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="426" swimtime="00:02:15.54" resultid="8511" heatid="10671" lane="7" entrytime="00:02:14.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                    <SPLIT distance="100" swimtime="00:01:05.49" />
                    <SPLIT distance="150" swimtime="00:01:40.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13068" nation="BRA" region="PR" clubid="8869" swrid="93787" name="Sociedade Morgenau" shortname="Morgenau">
          <ATHLETES>
            <ATHLETE firstname="Marcus" lastname="Vinicius De Almeida" birthdate="2009-06-16" gender="M" nation="BRA" license="348099" swrid="5600272" athleteid="8912" externalid="348099">
              <RESULTS>
                <RESULT eventid="1087" points="562" swimtime="00:02:32.02" resultid="8913" heatid="10492" lane="2" entrytime="00:02:34.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                    <SPLIT distance="100" swimtime="00:01:12.30" />
                    <SPLIT distance="150" swimtime="00:01:53.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="577" swimtime="00:00:31.16" resultid="8914" heatid="10575" lane="9" entrytime="00:00:31.76" entrycourse="LCM" />
                <RESULT eventid="1219" points="591" swimtime="00:01:07.76" resultid="8915" heatid="10599" lane="9" entrytime="00:01:08.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="478" swimtime="00:00:30.10" resultid="8916" heatid="10687" lane="0" entrytime="00:00:30.31" entrycourse="LCM" />
                <RESULT eventid="1273" points="473" swimtime="00:02:26.29" resultid="8917" heatid="10651" lane="2" entrytime="00:02:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                    <SPLIT distance="100" swimtime="00:01:12.98" />
                    <SPLIT distance="150" swimtime="00:01:51.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="452" swimtime="00:01:07.23" resultid="8918" heatid="10741" lane="4" entrytime="00:01:04.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Galarda" birthdate="2010-03-18" gender="M" nation="BRA" license="421438" swrid="5811239" athleteid="9024" externalid="421438">
              <RESULTS>
                <RESULT eventid="1103" points="282" swimtime="00:00:33.96" resultid="9025" heatid="10504" lane="8" entrytime="00:00:34.15" entrycourse="LCM" />
                <RESULT eventid="1187" points="160" swimtime="00:00:47.74" resultid="9026" heatid="10567" lane="4" />
                <RESULT eventid="1155" points="252" swimtime="00:01:13.39" resultid="9027" heatid="10535" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="290" swimtime="00:00:31.57" resultid="9028" heatid="10615" lane="4" entrytime="00:00:32.39" entrycourse="LCM" />
                <RESULT eventid="1305" points="185" swimtime="00:00:41.32" resultid="9029" heatid="10681" lane="4" />
                <RESULT eventid="1341" points="182" swimtime="00:01:27.14" resultid="9030" heatid="10703" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Gabriel Sarmento Buski" birthdate="2010-04-05" gender="M" nation="BRA" license="399533" swrid="5717264" athleteid="8933" externalid="399533">
              <RESULTS>
                <RESULT eventid="1123" points="449" swimtime="00:09:50.08" resultid="8934" heatid="10515" lane="2" entrytime="00:10:22.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                    <SPLIT distance="100" swimtime="00:01:07.15" />
                    <SPLIT distance="150" swimtime="00:01:44.01" />
                    <SPLIT distance="200" swimtime="00:02:19.95" />
                    <SPLIT distance="250" swimtime="00:02:57.58" />
                    <SPLIT distance="300" swimtime="00:03:34.71" />
                    <SPLIT distance="350" swimtime="00:04:12.86" />
                    <SPLIT distance="400" swimtime="00:04:49.95" />
                    <SPLIT distance="450" swimtime="00:05:28.09" />
                    <SPLIT distance="500" swimtime="00:06:05.69" />
                    <SPLIT distance="550" swimtime="00:06:44.47" />
                    <SPLIT distance="600" swimtime="00:07:23.09" />
                    <SPLIT distance="650" swimtime="00:08:00.43" />
                    <SPLIT distance="700" swimtime="00:08:38.17" />
                    <SPLIT distance="750" swimtime="00:09:15.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="373" swimtime="00:02:54.24" resultid="8935" heatid="10490" lane="7" entrytime="00:02:56.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.01" />
                    <SPLIT distance="100" swimtime="00:01:21.45" />
                    <SPLIT distance="150" swimtime="00:02:09.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="381" swimtime="00:00:35.79" resultid="8936" heatid="10572" lane="3" entrytime="00:00:38.66" entrycourse="LCM" />
                <RESULT eventid="1257" points="472" swimtime="00:18:37.63" resultid="8937" heatid="10636" lane="5" entrytime="00:19:01.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.80" />
                    <SPLIT distance="100" swimtime="00:01:06.52" />
                    <SPLIT distance="150" swimtime="00:01:43.00" />
                    <SPLIT distance="200" swimtime="00:02:19.70" />
                    <SPLIT distance="250" swimtime="00:02:56.66" />
                    <SPLIT distance="300" swimtime="00:03:34.19" />
                    <SPLIT distance="350" swimtime="00:04:11.48" />
                    <SPLIT distance="400" swimtime="00:04:48.47" />
                    <SPLIT distance="450" swimtime="00:05:27.25" />
                    <SPLIT distance="500" swimtime="00:06:04.85" />
                    <SPLIT distance="550" swimtime="00:06:43.24" />
                    <SPLIT distance="600" swimtime="00:07:21.04" />
                    <SPLIT distance="650" swimtime="00:07:59.75" />
                    <SPLIT distance="700" swimtime="00:08:37.27" />
                    <SPLIT distance="750" swimtime="00:09:14.76" />
                    <SPLIT distance="800" swimtime="00:09:52.16" />
                    <SPLIT distance="850" swimtime="00:10:29.93" />
                    <SPLIT distance="900" swimtime="00:11:07.32" />
                    <SPLIT distance="950" swimtime="00:11:45.13" />
                    <SPLIT distance="1000" swimtime="00:12:22.79" />
                    <SPLIT distance="1050" swimtime="00:13:00.93" />
                    <SPLIT distance="1100" swimtime="00:13:38.40" />
                    <SPLIT distance="1150" swimtime="00:14:16.24" />
                    <SPLIT distance="1200" swimtime="00:14:54.64" />
                    <SPLIT distance="1250" swimtime="00:15:33.53" />
                    <SPLIT distance="1300" swimtime="00:16:11.05" />
                    <SPLIT distance="1350" swimtime="00:16:49.74" />
                    <SPLIT distance="1400" swimtime="00:17:26.90" />
                    <SPLIT distance="1450" swimtime="00:18:03.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="373" swimtime="00:01:18.99" resultid="8938" heatid="10596" lane="4" entrytime="00:01:18.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="457" swimtime="00:04:45.67" resultid="8939" heatid="10721" lane="5" entrytime="00:04:53.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                    <SPLIT distance="100" swimtime="00:01:04.15" />
                    <SPLIT distance="150" swimtime="00:01:40.13" />
                    <SPLIT distance="200" swimtime="00:02:16.51" />
                    <SPLIT distance="250" swimtime="00:02:53.84" />
                    <SPLIT distance="300" swimtime="00:03:31.67" />
                    <SPLIT distance="350" swimtime="00:04:09.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Riccieri" lastname="Rodrigues Muzolon" birthdate="2010-11-08" gender="M" nation="BRA" license="385439" swrid="5588887" athleteid="8945" externalid="385439">
              <RESULTS>
                <RESULT eventid="1123" points="364" swimtime="00:10:32.83" resultid="8946" heatid="10517" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                    <SPLIT distance="100" swimtime="00:01:09.56" />
                    <SPLIT distance="150" swimtime="00:01:47.33" />
                    <SPLIT distance="200" swimtime="00:02:26.37" />
                    <SPLIT distance="250" swimtime="00:03:06.31" />
                    <SPLIT distance="300" swimtime="00:03:46.74" />
                    <SPLIT distance="350" swimtime="00:04:27.50" />
                    <SPLIT distance="400" swimtime="00:05:08.42" />
                    <SPLIT distance="450" swimtime="00:05:50.10" />
                    <SPLIT distance="500" swimtime="00:06:30.84" />
                    <SPLIT distance="550" swimtime="00:07:11.54" />
                    <SPLIT distance="600" swimtime="00:07:52.59" />
                    <SPLIT distance="650" swimtime="00:08:33.13" />
                    <SPLIT distance="700" swimtime="00:09:13.71" />
                    <SPLIT distance="750" swimtime="00:09:53.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="351" swimtime="00:20:33.78" resultid="8947" heatid="10637" lane="7" entrytime="00:20:37.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.87" />
                    <SPLIT distance="100" swimtime="00:01:11.29" />
                    <SPLIT distance="150" swimtime="00:01:49.68" />
                    <SPLIT distance="200" swimtime="00:02:29.36" />
                    <SPLIT distance="250" swimtime="00:03:09.20" />
                    <SPLIT distance="300" swimtime="00:03:49.28" />
                    <SPLIT distance="350" swimtime="00:04:30.05" />
                    <SPLIT distance="400" swimtime="00:05:11.43" />
                    <SPLIT distance="450" swimtime="00:05:53.60" />
                    <SPLIT distance="500" swimtime="00:06:35.11" />
                    <SPLIT distance="550" swimtime="00:07:17.05" />
                    <SPLIT distance="600" swimtime="00:07:59.28" />
                    <SPLIT distance="650" swimtime="00:08:41.32" />
                    <SPLIT distance="700" swimtime="00:09:22.78" />
                    <SPLIT distance="750" swimtime="00:10:05.01" />
                    <SPLIT distance="800" swimtime="00:10:47.40" />
                    <SPLIT distance="850" swimtime="00:11:29.59" />
                    <SPLIT distance="900" swimtime="00:12:11.02" />
                    <SPLIT distance="950" swimtime="00:12:52.65" />
                    <SPLIT distance="1000" swimtime="00:13:34.93" />
                    <SPLIT distance="1050" swimtime="00:14:17.06" />
                    <SPLIT distance="1100" swimtime="00:14:58.88" />
                    <SPLIT distance="1150" swimtime="00:15:41.75" />
                    <SPLIT distance="1200" swimtime="00:16:23.87" />
                    <SPLIT distance="1250" swimtime="00:17:06.23" />
                    <SPLIT distance="1300" swimtime="00:17:48.46" />
                    <SPLIT distance="1350" swimtime="00:18:30.10" />
                    <SPLIT distance="1400" swimtime="00:19:11.98" />
                    <SPLIT distance="1450" swimtime="00:19:53.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="321" swimtime="00:01:23.04" resultid="8948" heatid="10594" lane="5" entrytime="00:01:26.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="389" swimtime="00:02:19.61" resultid="8949" heatid="10666" lane="3" entrytime="00:02:34.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                    <SPLIT distance="100" swimtime="00:01:07.99" />
                    <SPLIT distance="150" swimtime="00:01:43.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="358" swimtime="00:01:12.65" resultid="8950" heatid="10737" lane="4" entrytime="00:01:16.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabryel" lastname="Denk" birthdate="2011-05-09" gender="M" nation="BRA" license="391138" swrid="5602531" athleteid="8970" externalid="391138">
              <RESULTS>
                <RESULT eventid="1123" points="425" swimtime="00:10:01.12" resultid="8971" heatid="10515" lane="8" entrytime="00:10:26.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                    <SPLIT distance="100" swimtime="00:01:06.85" />
                    <SPLIT distance="150" swimtime="00:01:43.71" />
                    <SPLIT distance="200" swimtime="00:02:21.36" />
                    <SPLIT distance="250" swimtime="00:02:59.64" />
                    <SPLIT distance="300" swimtime="00:03:38.14" />
                    <SPLIT distance="350" swimtime="00:04:17.43" />
                    <SPLIT distance="400" swimtime="00:04:56.89" />
                    <SPLIT distance="450" swimtime="00:05:35.55" />
                    <SPLIT distance="500" swimtime="00:06:14.26" />
                    <SPLIT distance="550" swimtime="00:06:53.21" />
                    <SPLIT distance="600" swimtime="00:07:31.17" />
                    <SPLIT distance="650" swimtime="00:08:09.65" />
                    <SPLIT distance="700" swimtime="00:08:47.98" />
                    <SPLIT distance="750" swimtime="00:09:26.06" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 6.4 - Não começou a executar a virada imediatamente após virar para a posição de peito.  (Horário: 9:41), Na volta dos 50 e 150m." eventid="1071" status="DSQ" swimtime="00:02:37.31" resultid="8972" heatid="10477" lane="8" entrytime="00:02:44.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.83" />
                    <SPLIT distance="100" swimtime="00:01:16.70" />
                    <SPLIT distance="150" swimtime="00:01:58.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="359" swimtime="00:01:05.24" resultid="8973" heatid="10544" lane="2" entrytime="00:01:06.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="440" swimtime="00:19:04.03" resultid="8974" heatid="10636" lane="3" entrytime="00:19:01.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.87" />
                    <SPLIT distance="100" swimtime="00:01:07.06" />
                    <SPLIT distance="150" swimtime="00:01:44.69" />
                    <SPLIT distance="200" swimtime="00:02:22.07" />
                    <SPLIT distance="250" swimtime="00:02:59.52" />
                    <SPLIT distance="300" swimtime="00:03:37.92" />
                    <SPLIT distance="350" swimtime="00:04:15.39" />
                    <SPLIT distance="400" swimtime="00:04:53.46" />
                    <SPLIT distance="450" swimtime="00:05:31.37" />
                    <SPLIT distance="500" swimtime="00:06:09.74" />
                    <SPLIT distance="550" swimtime="00:06:48.03" />
                    <SPLIT distance="600" swimtime="00:07:26.25" />
                    <SPLIT distance="650" swimtime="00:08:04.89" />
                    <SPLIT distance="700" swimtime="00:08:43.39" />
                    <SPLIT distance="750" swimtime="00:09:21.69" />
                    <SPLIT distance="800" swimtime="00:10:00.56" />
                    <SPLIT distance="850" swimtime="00:10:39.18" />
                    <SPLIT distance="900" swimtime="00:11:17.89" />
                    <SPLIT distance="950" swimtime="00:11:56.53" />
                    <SPLIT distance="1000" swimtime="00:12:35.60" />
                    <SPLIT distance="1050" swimtime="00:13:14.40" />
                    <SPLIT distance="1100" swimtime="00:13:53.11" />
                    <SPLIT distance="1150" swimtime="00:14:32.02" />
                    <SPLIT distance="1200" swimtime="00:15:11.48" />
                    <SPLIT distance="1250" swimtime="00:15:50.09" />
                    <SPLIT distance="1300" swimtime="00:16:29.71" />
                    <SPLIT distance="1350" swimtime="00:17:08.48" />
                    <SPLIT distance="1400" swimtime="00:17:48.29" />
                    <SPLIT distance="1450" swimtime="00:18:26.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="419" swimtime="00:04:53.88" resultid="8975" heatid="10721" lane="6" entrytime="00:04:54.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                    <SPLIT distance="100" swimtime="00:01:07.08" />
                    <SPLIT distance="150" swimtime="00:01:44.67" />
                    <SPLIT distance="200" swimtime="00:02:22.78" />
                    <SPLIT distance="250" swimtime="00:03:01.45" />
                    <SPLIT distance="300" swimtime="00:03:39.77" />
                    <SPLIT distance="350" swimtime="00:04:17.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="324" swimtime="00:01:15.11" resultid="8976" heatid="10738" lane="7" entrytime="00:01:14.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luana" lastname="Yoshie Kimura" birthdate="2010-07-08" gender="F" nation="BRA" license="391142" swrid="5600277" athleteid="8870" externalid="391142">
              <RESULTS>
                <RESULT eventid="1079" points="477" swimtime="00:02:56.03" resultid="8871" heatid="10485" lane="6" entrytime="00:02:57.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.65" />
                    <SPLIT distance="100" swimtime="00:01:20.85" />
                    <SPLIT distance="150" swimtime="00:02:08.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="502" swimtime="00:00:36.69" resultid="8872" heatid="10565" lane="2" entrytime="00:00:36.06" entrycourse="LCM" />
                <RESULT eventid="1131" points="373" swimtime="00:06:06.97" resultid="8873" heatid="10520" lane="9" entrytime="00:06:05.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                    <SPLIT distance="100" swimtime="00:01:23.35" />
                    <SPLIT distance="150" swimtime="00:02:13.79" />
                    <SPLIT distance="200" swimtime="00:03:04.10" />
                    <SPLIT distance="250" swimtime="00:03:51.38" />
                    <SPLIT distance="300" swimtime="00:04:39.66" />
                    <SPLIT distance="350" swimtime="00:05:25.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="356" swimtime="00:11:23.85" resultid="8874" heatid="10633" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                    <SPLIT distance="100" swimtime="00:01:16.08" />
                    <SPLIT distance="150" swimtime="00:01:58.01" />
                    <SPLIT distance="200" swimtime="00:02:40.53" />
                    <SPLIT distance="250" swimtime="00:03:23.53" />
                    <SPLIT distance="300" swimtime="00:04:06.92" />
                    <SPLIT distance="350" swimtime="00:04:51.80" />
                    <SPLIT distance="400" swimtime="00:05:35.83" />
                    <SPLIT distance="450" swimtime="00:06:20.07" />
                    <SPLIT distance="500" swimtime="00:07:04.06" />
                    <SPLIT distance="550" swimtime="00:07:48.30" />
                    <SPLIT distance="600" swimtime="00:08:32.36" />
                    <SPLIT distance="650" swimtime="00:09:16.91" />
                    <SPLIT distance="700" swimtime="00:10:00.57" />
                    <SPLIT distance="750" swimtime="00:10:42.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="511" swimtime="00:01:20.20" resultid="8875" heatid="10589" lane="8" entrytime="00:01:19.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="399" swimtime="00:02:51.20" resultid="8876" heatid="10643" lane="9" entrytime="00:02:47.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                    <SPLIT distance="100" swimtime="00:01:25.54" />
                    <SPLIT distance="150" swimtime="00:02:11.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Capoia Soares" birthdate="2011-11-07" gender="M" nation="BRA" license="393257" swrid="5616440" athleteid="8991" externalid="393257">
              <RESULTS>
                <RESULT eventid="1103" points="159" swimtime="00:00:41.07" resultid="8992" heatid="10502" lane="3" entrytime="00:00:55.50" entrycourse="LCM" />
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 18:53), 150m" eventid="1171" status="DSQ" swimtime="00:03:20.74" resultid="8993" heatid="10555" lane="5" entrytime="00:03:22.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.07" />
                    <SPLIT distance="100" swimtime="00:01:32.37" />
                    <SPLIT distance="150" swimtime="00:02:27.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="217" swimtime="00:00:34.76" resultid="8994" heatid="10612" lane="4" />
                <RESULT eventid="1341" points="161" swimtime="00:01:30.80" resultid="8995" heatid="10705" lane="8" entrytime="00:01:33.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanne" lastname="Gomes" birthdate="2008-03-20" gender="M" nation="BRA" license="421442" swrid="5768391" athleteid="9051" externalid="421442">
              <RESULTS>
                <RESULT eventid="1103" points="260" swimtime="00:00:34.88" resultid="9052" heatid="10499" lane="4" />
                <RESULT eventid="1087" points="360" swimtime="00:02:56.27" resultid="9053" heatid="10490" lane="8" entrytime="00:02:57.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.13" />
                    <SPLIT distance="100" swimtime="00:01:22.54" />
                    <SPLIT distance="150" swimtime="00:02:10.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="326" swimtime="00:00:37.68" resultid="9054" heatid="10573" lane="0" entrytime="00:00:36.54" entrycourse="LCM" />
                <RESULT eventid="1155" points="328" swimtime="00:01:07.28" resultid="9055" heatid="10536" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="326" swimtime="00:01:22.59" resultid="9056" heatid="10596" lane="3" entrytime="00:01:18.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="338" swimtime="00:02:26.38" resultid="9057" heatid="10661" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                    <SPLIT distance="100" swimtime="00:01:08.64" />
                    <SPLIT distance="150" swimtime="00:01:47.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Rafaella Dos Santos" birthdate="2005-02-25" gender="F" nation="BRA" license="358849" swrid="5757094" athleteid="8877" externalid="358849">
              <RESULTS>
                <RESULT eventid="1079" points="288" swimtime="00:03:28.14" resultid="8878" heatid="10482" lane="5" entrytime="00:03:20.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.03" />
                    <SPLIT distance="100" swimtime="00:01:35.16" />
                    <SPLIT distance="150" swimtime="00:02:32.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="330" swimtime="00:00:42.17" resultid="8879" heatid="10563" lane="8" entrytime="00:00:41.85" entrycourse="LCM" />
                <RESULT eventid="1211" points="309" swimtime="00:01:34.76" resultid="8880" heatid="10585" lane="6" entrytime="00:01:31.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="273" swimtime="00:03:14.38" resultid="8881" heatid="10640" lane="7" entrytime="00:03:15.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.49" />
                    <SPLIT distance="100" swimtime="00:01:35.79" />
                    <SPLIT distance="150" swimtime="00:02:30.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="258" swimtime="00:02:56.29" resultid="8882" heatid="10654" lane="6" entrytime="00:02:56.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.62" />
                    <SPLIT distance="100" swimtime="00:01:24.82" />
                    <SPLIT distance="150" swimtime="00:02:12.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Clara Martins" birthdate="2012-12-03" gender="F" nation="BRA" license="421441" swrid="5505965" athleteid="9044" externalid="421441">
              <RESULTS>
                <RESULT eventid="1095" points="185" swimtime="00:00:42.82" resultid="9045" heatid="10493" lane="3" />
                <RESULT eventid="1079" points="266" swimtime="00:03:33.87" resultid="9046" heatid="10482" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.09" />
                    <SPLIT distance="100" swimtime="00:01:40.55" />
                    <SPLIT distance="150" swimtime="00:02:37.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="335" swimtime="00:01:14.39" resultid="9047" heatid="10525" lane="9" />
                <RESULT eventid="1249" points="344" swimtime="00:11:31.38" resultid="9048" heatid="10633" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                    <SPLIT distance="100" swimtime="00:01:16.56" />
                    <SPLIT distance="150" swimtime="00:01:58.94" />
                    <SPLIT distance="200" swimtime="00:02:43.04" />
                    <SPLIT distance="250" swimtime="00:03:27.44" />
                    <SPLIT distance="300" swimtime="00:04:11.48" />
                    <SPLIT distance="350" swimtime="00:04:55.41" />
                    <SPLIT distance="400" swimtime="00:05:39.59" />
                    <SPLIT distance="450" swimtime="00:06:23.74" />
                    <SPLIT distance="500" swimtime="00:07:07.94" />
                    <SPLIT distance="550" swimtime="00:07:52.22" />
                    <SPLIT distance="600" swimtime="00:08:36.96" />
                    <SPLIT distance="650" swimtime="00:09:20.98" />
                    <SPLIT distance="700" swimtime="00:10:02.84" />
                    <SPLIT distance="750" swimtime="00:10:46.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="290" swimtime="00:01:36.88" resultid="9049" heatid="10584" lane="7" entrytime="00:01:39.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="353" swimtime="00:05:32.80" resultid="9050" heatid="10713" lane="4" entrytime="00:05:30.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                    <SPLIT distance="100" swimtime="00:01:16.29" />
                    <SPLIT distance="150" swimtime="00:01:59.17" />
                    <SPLIT distance="200" swimtime="00:02:42.12" />
                    <SPLIT distance="250" swimtime="00:03:25.05" />
                    <SPLIT distance="300" swimtime="00:04:08.62" />
                    <SPLIT distance="350" swimtime="00:04:51.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Andreis Ramos" birthdate="2007-03-26" gender="M" nation="BRA" license="406719" swrid="5717243" athleteid="8940" externalid="406719">
              <RESULTS>
                <RESULT eventid="1103" points="316" swimtime="00:00:32.69" resultid="8941" heatid="10505" lane="3" entrytime="00:00:31.35" entrycourse="LCM" />
                <RESULT eventid="1155" points="414" swimtime="00:01:02.25" resultid="8942" heatid="10548" lane="9" entrytime="00:01:01.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="365" swimtime="00:02:22.70" resultid="8943" heatid="10668" lane="8" entrytime="00:02:23.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                    <SPLIT distance="100" swimtime="00:01:07.87" />
                    <SPLIT distance="150" swimtime="00:01:45.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="386" swimtime="00:05:02.22" resultid="8944" heatid="10720" lane="9" entrytime="00:05:16.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                    <SPLIT distance="100" swimtime="00:01:10.01" />
                    <SPLIT distance="150" swimtime="00:01:49.71" />
                    <SPLIT distance="200" swimtime="00:02:29.32" />
                    <SPLIT distance="250" swimtime="00:03:09.58" />
                    <SPLIT distance="300" swimtime="00:03:48.35" />
                    <SPLIT distance="350" swimtime="00:04:27.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Geovana" lastname="Dos Santos" birthdate="2011-01-20" gender="F" nation="BRA" license="367254" swrid="5602533" athleteid="8883" externalid="367254">
              <RESULTS>
                <RESULT eventid="1063" points="307" swimtime="00:03:02.53" resultid="8884" heatid="10470" lane="6" entrytime="00:03:02.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="325" swimtime="00:01:15.19" resultid="8885" heatid="10527" lane="7" entrytime="00:01:15.96" entrycourse="LCM" />
                <RESULT eventid="1297" points="314" swimtime="00:00:39.51" resultid="8886" heatid="10679" lane="8" entrytime="00:00:39.25" entrycourse="LCM" />
                <RESULT eventid="1281" points="323" swimtime="00:02:43.57" resultid="8887" heatid="10655" lane="2" entrytime="00:02:39.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.92" />
                    <SPLIT distance="100" swimtime="00:01:18.02" />
                    <SPLIT distance="150" swimtime="00:02:01.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="313" swimtime="00:05:46.66" resultid="8888" heatid="10713" lane="8" entrytime="00:05:46.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.43" />
                    <SPLIT distance="100" swimtime="00:01:19.62" />
                    <SPLIT distance="150" swimtime="00:02:04.14" />
                    <SPLIT distance="200" swimtime="00:02:48.84" />
                    <SPLIT distance="250" swimtime="00:03:34.33" />
                    <SPLIT distance="300" swimtime="00:04:18.55" />
                    <SPLIT distance="350" swimtime="00:05:04.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="282" swimtime="00:01:27.04" resultid="8889" heatid="10729" lane="9" entrytime="00:01:24.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hayanna" lastname="Piovezan" birthdate="1996-06-25" gender="F" nation="BRA" license="100002" athleteid="8895" externalid="100002">
              <RESULTS>
                <RESULT eventid="1179" points="392" swimtime="00:00:39.82" resultid="8896" heatid="10561" lane="7" />
                <RESULT eventid="1211" points="341" swimtime="00:01:31.79" resultid="8897" heatid="10583" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Henrique Opuchkevich" birthdate="2011-02-22" gender="M" nation="BRA" license="406720" swrid="5717273" athleteid="9003" externalid="406720">
              <RESULTS>
                <RESULT eventid="1123" points="391" swimtime="00:10:18.04" resultid="9004" heatid="10515" lane="0" entrytime="00:10:27.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                    <SPLIT distance="100" swimtime="00:01:10.70" />
                    <SPLIT distance="150" swimtime="00:01:50.10" />
                    <SPLIT distance="200" swimtime="00:02:29.07" />
                    <SPLIT distance="250" swimtime="00:03:08.92" />
                    <SPLIT distance="300" swimtime="00:03:48.43" />
                    <SPLIT distance="350" swimtime="00:04:28.51" />
                    <SPLIT distance="400" swimtime="00:05:08.20" />
                    <SPLIT distance="450" swimtime="00:05:48.02" />
                    <SPLIT distance="500" swimtime="00:06:27.83" />
                    <SPLIT distance="550" swimtime="00:07:07.40" />
                    <SPLIT distance="600" swimtime="00:07:47.00" />
                    <SPLIT distance="650" swimtime="00:08:27.13" />
                    <SPLIT distance="700" swimtime="00:09:05.09" />
                    <SPLIT distance="750" swimtime="00:09:42.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="380" swimtime="00:02:53.12" resultid="9005" heatid="10491" lane="9" entrytime="00:02:52.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.37" />
                    <SPLIT distance="100" swimtime="00:01:21.22" />
                    <SPLIT distance="150" swimtime="00:02:07.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="368" swimtime="00:00:36.21" resultid="9006" heatid="10572" lane="4" entrytime="00:00:37.02" entrycourse="LCM" />
                <RESULT eventid="1257" points="433" swimtime="00:19:10.83" resultid="9007" heatid="10636" lane="0" entrytime="00:19:33.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                    <SPLIT distance="100" swimtime="00:01:09.03" />
                    <SPLIT distance="150" swimtime="00:01:48.20" />
                    <SPLIT distance="200" swimtime="00:02:26.75" />
                    <SPLIT distance="250" swimtime="00:03:06.31" />
                    <SPLIT distance="300" swimtime="00:03:45.42" />
                    <SPLIT distance="350" swimtime="00:04:25.06" />
                    <SPLIT distance="400" swimtime="00:05:03.91" />
                    <SPLIT distance="450" swimtime="00:05:43.13" />
                    <SPLIT distance="500" swimtime="00:06:21.91" />
                    <SPLIT distance="550" swimtime="00:07:00.98" />
                    <SPLIT distance="600" swimtime="00:07:39.88" />
                    <SPLIT distance="650" swimtime="00:08:18.58" />
                    <SPLIT distance="700" swimtime="00:08:57.09" />
                    <SPLIT distance="750" swimtime="00:09:35.54" />
                    <SPLIT distance="800" swimtime="00:10:13.87" />
                    <SPLIT distance="850" swimtime="00:10:52.69" />
                    <SPLIT distance="900" swimtime="00:11:31.78" />
                    <SPLIT distance="950" swimtime="00:12:10.57" />
                    <SPLIT distance="1000" swimtime="00:12:48.11" />
                    <SPLIT distance="1050" swimtime="00:13:27.03" />
                    <SPLIT distance="1100" swimtime="00:14:05.16" />
                    <SPLIT distance="1150" swimtime="00:14:44.47" />
                    <SPLIT distance="1200" swimtime="00:15:23.00" />
                    <SPLIT distance="1250" swimtime="00:16:01.71" />
                    <SPLIT distance="1300" swimtime="00:16:40.73" />
                    <SPLIT distance="1350" swimtime="00:17:19.88" />
                    <SPLIT distance="1400" swimtime="00:17:57.79" />
                    <SPLIT distance="1450" swimtime="00:18:35.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="342" swimtime="00:01:21.26" resultid="9008" heatid="10596" lane="1" entrytime="00:01:20.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="329" swimtime="00:02:45.12" resultid="9009" heatid="10649" lane="9" entrytime="00:02:44.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                    <SPLIT distance="100" swimtime="00:01:23.41" />
                    <SPLIT distance="150" swimtime="00:02:07.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Tomaz Zmievski" birthdate="2012-09-20" gender="F" nation="BRA" license="406725" swrid="5717300" athleteid="9017" externalid="406725">
              <RESULTS>
                <RESULT eventid="1115" points="275" swimtime="00:23:34.78" resultid="9018" heatid="10512" lane="9">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                    <SPLIT distance="100" swimtime="00:01:25.47" />
                    <SPLIT distance="150" swimtime="00:02:13.14" />
                    <SPLIT distance="200" swimtime="00:03:01.32" />
                    <SPLIT distance="250" swimtime="00:03:47.27" />
                    <SPLIT distance="300" swimtime="00:04:34.30" />
                    <SPLIT distance="350" swimtime="00:05:22.70" />
                    <SPLIT distance="400" swimtime="00:06:10.33" />
                    <SPLIT distance="450" swimtime="00:06:57.03" />
                    <SPLIT distance="500" swimtime="00:07:45.31" />
                    <SPLIT distance="550" swimtime="00:08:34.83" />
                    <SPLIT distance="600" swimtime="00:09:22.85" />
                    <SPLIT distance="650" swimtime="00:10:11.40" />
                    <SPLIT distance="700" swimtime="00:10:58.80" />
                    <SPLIT distance="750" swimtime="00:11:45.28" />
                    <SPLIT distance="800" swimtime="00:12:33.08" />
                    <SPLIT distance="850" swimtime="00:13:21.48" />
                    <SPLIT distance="900" swimtime="00:14:08.88" />
                    <SPLIT distance="950" swimtime="00:14:56.91" />
                    <SPLIT distance="1000" swimtime="00:15:44.67" />
                    <SPLIT distance="1050" swimtime="00:16:32.23" />
                    <SPLIT distance="1100" swimtime="00:17:20.95" />
                    <SPLIT distance="1150" swimtime="00:18:08.98" />
                    <SPLIT distance="1200" swimtime="00:18:56.68" />
                    <SPLIT distance="1250" swimtime="00:19:43.45" />
                    <SPLIT distance="1300" swimtime="00:20:30.60" />
                    <SPLIT distance="1350" swimtime="00:21:18.60" />
                    <SPLIT distance="1400" swimtime="00:22:06.33" />
                    <SPLIT distance="1450" swimtime="00:22:52.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="320" swimtime="00:01:15.54" resultid="9019" heatid="10526" lane="1" entrytime="00:01:20.53" entrycourse="LCM" />
                <RESULT eventid="1249" points="300" swimtime="00:12:04.10" resultid="9020" heatid="10634" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.82" />
                    <SPLIT distance="100" swimtime="00:01:20.76" />
                    <SPLIT distance="150" swimtime="00:02:06.61" />
                    <SPLIT distance="200" swimtime="00:02:52.37" />
                    <SPLIT distance="250" swimtime="00:03:38.57" />
                    <SPLIT distance="300" swimtime="00:04:25.11" />
                    <SPLIT distance="350" swimtime="00:05:12.26" />
                    <SPLIT distance="400" swimtime="00:05:58.55" />
                    <SPLIT distance="450" swimtime="00:06:45.35" />
                    <SPLIT distance="500" swimtime="00:07:31.67" />
                    <SPLIT distance="550" swimtime="00:08:18.34" />
                    <SPLIT distance="600" swimtime="00:09:04.12" />
                    <SPLIT distance="650" swimtime="00:09:49.72" />
                    <SPLIT distance="700" swimtime="00:10:35.25" />
                    <SPLIT distance="750" swimtime="00:11:20.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="260" swimtime="00:03:17.60" resultid="9021" heatid="10640" lane="1" entrytime="00:03:16.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.02" />
                    <SPLIT distance="100" swimtime="00:01:36.40" />
                    <SPLIT distance="150" swimtime="00:02:36.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="294" swimtime="00:02:48.60" resultid="9022" heatid="10654" lane="3" entrytime="00:02:54.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                    <SPLIT distance="100" swimtime="00:01:20.68" />
                    <SPLIT distance="150" swimtime="00:02:05.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="301" swimtime="00:05:50.90" resultid="9023" heatid="10712" lane="5" entrytime="00:06:04.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                    <SPLIT distance="100" swimtime="00:01:20.78" />
                    <SPLIT distance="150" swimtime="00:02:05.86" />
                    <SPLIT distance="200" swimtime="00:02:51.63" />
                    <SPLIT distance="250" swimtime="00:03:37.29" />
                    <SPLIT distance="300" swimtime="00:04:22.68" />
                    <SPLIT distance="350" swimtime="00:05:07.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Eduardo Gavinski Alves" birthdate="2012-10-12" gender="M" nation="BRA" license="369324" swrid="5588674" athleteid="8951" externalid="369324">
              <RESULTS>
                <RESULT eventid="1071" points="302" swimtime="00:02:46.72" resultid="8952" heatid="10476" lane="5" entrytime="00:02:45.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.82" />
                    <SPLIT distance="100" swimtime="00:01:22.92" />
                    <SPLIT distance="150" swimtime="00:02:05.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="294" swimtime="00:01:09.72" resultid="8953" heatid="10542" lane="9" entrytime="00:01:10.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="303" swimtime="00:00:31.10" resultid="8954" heatid="10616" lane="6" entrytime="00:00:32.01" entrycourse="LCM" />
                <RESULT eventid="1305" points="303" swimtime="00:00:35.06" resultid="8955" heatid="10685" lane="6" entrytime="00:00:34.93" entrycourse="LCM" />
                <RESULT eventid="1273" points="277" swimtime="00:02:54.81" resultid="8956" heatid="10647" lane="4" entrytime="00:02:55.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.76" />
                    <SPLIT distance="100" swimtime="00:01:23.12" />
                    <SPLIT distance="150" swimtime="00:02:17.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1373" points="288" swimtime="00:01:18.13" resultid="8957" heatid="10738" lane="9" entrytime="00:01:15.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Liz Skowronski" birthdate="2008-01-24" gender="F" nation="BRA" license="358245" swrid="5600202" athleteid="8898" externalid="358245">
              <RESULTS>
                <RESULT eventid="1115" points="349" swimtime="00:21:46.70" resultid="8899" heatid="10512" lane="7" entrytime="00:21:17.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.19" />
                    <SPLIT distance="100" swimtime="00:01:19.84" />
                    <SPLIT distance="150" swimtime="00:02:02.84" />
                    <SPLIT distance="200" swimtime="00:02:45.52" />
                    <SPLIT distance="250" swimtime="00:03:28.93" />
                    <SPLIT distance="300" swimtime="00:04:12.55" />
                    <SPLIT distance="350" swimtime="00:04:56.48" />
                    <SPLIT distance="400" swimtime="00:05:40.06" />
                    <SPLIT distance="450" swimtime="00:06:24.00" />
                    <SPLIT distance="500" swimtime="00:07:07.58" />
                    <SPLIT distance="550" swimtime="00:07:51.67" />
                    <SPLIT distance="600" swimtime="00:08:34.88" />
                    <SPLIT distance="650" swimtime="00:09:18.69" />
                    <SPLIT distance="700" swimtime="00:10:02.68" />
                    <SPLIT distance="750" swimtime="00:10:47.17" />
                    <SPLIT distance="800" swimtime="00:11:31.27" />
                    <SPLIT distance="850" swimtime="00:12:16.02" />
                    <SPLIT distance="900" swimtime="00:12:59.70" />
                    <SPLIT distance="950" swimtime="00:13:44.73" />
                    <SPLIT distance="1000" swimtime="00:14:29.00" />
                    <SPLIT distance="1050" swimtime="00:15:13.95" />
                    <SPLIT distance="1100" swimtime="00:15:57.86" />
                    <SPLIT distance="1150" swimtime="00:16:42.47" />
                    <SPLIT distance="1200" swimtime="00:17:26.20" />
                    <SPLIT distance="1250" swimtime="00:18:10.18" />
                    <SPLIT distance="1300" swimtime="00:18:53.90" />
                    <SPLIT distance="1350" swimtime="00:19:37.82" />
                    <SPLIT distance="1400" swimtime="00:20:20.93" />
                    <SPLIT distance="1450" swimtime="00:21:04.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="260" swimtime="00:00:38.23" resultid="8900" heatid="10495" lane="9" />
                <RESULT eventid="1163" points="202" swimtime="00:03:27.30" resultid="8901" heatid="10553" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.24" />
                    <SPLIT distance="150" swimtime="00:02:29.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="311" swimtime="00:06:29.89" resultid="8902" heatid="10519" lane="0" entrytime="00:06:19.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                    <SPLIT distance="100" swimtime="00:01:27.81" />
                    <SPLIT distance="150" swimtime="00:02:18.39" />
                    <SPLIT distance="200" swimtime="00:03:07.77" />
                    <SPLIT distance="300" swimtime="00:05:02.60" />
                    <SPLIT distance="350" swimtime="00:05:47.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="329" swimtime="00:03:02.65" resultid="8903" heatid="10641" lane="4" entrytime="00:02:54.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                    <SPLIT distance="150" swimtime="00:02:20.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="249" swimtime="00:01:27.65" resultid="8904" heatid="10700" lane="1" entrytime="00:01:30.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Eduardo Hoinatski" birthdate="2011-12-30" gender="M" nation="BRA" license="423406" athleteid="9068" externalid="423406">
              <RESULTS>
                <RESULT eventid="1071" points="163" swimtime="00:03:24.72" resultid="9069" heatid="10474" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.30" />
                    <SPLIT distance="150" swimtime="00:02:33.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="129" swimtime="00:00:51.29" resultid="9070" heatid="10569" lane="0" />
                <RESULT eventid="1155" points="224" swimtime="00:01:16.31" resultid="9071" heatid="10536" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="216" swimtime="00:00:34.80" resultid="9072" heatid="10611" lane="0" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabella" lastname="Denez" birthdate="2011-04-25" gender="F" nation="BRA" license="421439" swrid="5775839" athleteid="9031" externalid="421439">
              <RESULTS>
                <RESULT eventid="1095" points="178" swimtime="00:00:43.35" resultid="9032" heatid="10493" lane="4" />
                <RESULT eventid="1147" points="242" swimtime="00:01:22.89" resultid="9033" heatid="10525" lane="2" entrytime="00:01:23.36" entrycourse="LCM" />
                <RESULT eventid="1211" points="203" swimtime="00:01:49.10" resultid="9034" heatid="10584" lane="9" entrytime="00:01:43.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="235" swimtime="00:00:43.47" resultid="9035" heatid="10676" lane="8" />
                <RESULT eventid="1281" points="271" swimtime="00:02:53.26" resultid="9036" heatid="10654" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.57" />
                    <SPLIT distance="100" swimtime="00:01:24.46" />
                    <SPLIT distance="150" swimtime="00:02:10.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="232" swimtime="00:01:32.85" resultid="9037" heatid="10727" lane="2" entrytime="00:01:34.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolas" lastname="Mingorance Martins" birthdate="2007-10-13" gender="M" nation="BRA" license="393920" swrid="5622295" athleteid="8919" externalid="393920">
              <RESULTS>
                <RESULT eventid="1071" points="394" swimtime="00:02:32.58" resultid="8920" heatid="10478" lane="9" entrytime="00:02:34.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                    <SPLIT distance="100" swimtime="00:01:12.49" />
                    <SPLIT distance="150" swimtime="00:01:52.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="560" swimtime="00:00:56.26" resultid="8921" heatid="10551" lane="9" entrytime="00:00:56.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="540" swimtime="00:00:25.67" resultid="8922" heatid="10626" lane="3" entrytime="00:00:25.67" entrycourse="LCM" />
                <RESULT eventid="1305" points="411" swimtime="00:00:31.65" resultid="8923" heatid="10681" lane="9" />
                <RESULT eventid="1289" points="535" swimtime="00:02:05.59" resultid="8924" heatid="10673" lane="8" entrytime="00:02:06.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.12" />
                    <SPLIT distance="100" swimtime="00:00:59.42" />
                    <SPLIT distance="150" swimtime="00:01:32.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="480" swimtime="00:04:41.04" resultid="8925" heatid="10722" lane="2" entrytime="00:04:44.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                    <SPLIT distance="100" swimtime="00:01:05.07" />
                    <SPLIT distance="150" swimtime="00:01:40.07" />
                    <SPLIT distance="200" swimtime="00:02:15.48" />
                    <SPLIT distance="250" swimtime="00:02:51.53" />
                    <SPLIT distance="300" swimtime="00:03:28.26" />
                    <SPLIT distance="350" swimtime="00:04:04.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benito" lastname="Alves Sant&apos;Ana" birthdate="2009-06-01" gender="M" nation="BRA" license="376585" swrid="5351951" athleteid="8905" externalid="376585">
              <RESULTS>
                <RESULT eventid="1123" points="566" swimtime="00:09:06.36" resultid="8906" heatid="10513" lane="7" entrytime="00:09:08.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.58" />
                    <SPLIT distance="100" swimtime="00:01:01.85" />
                    <SPLIT distance="150" swimtime="00:01:35.34" />
                    <SPLIT distance="200" swimtime="00:02:09.41" />
                    <SPLIT distance="250" swimtime="00:02:43.92" />
                    <SPLIT distance="300" swimtime="00:03:18.27" />
                    <SPLIT distance="350" swimtime="00:03:53.42" />
                    <SPLIT distance="400" swimtime="00:04:28.36" />
                    <SPLIT distance="450" swimtime="00:05:03.71" />
                    <SPLIT distance="500" swimtime="00:05:38.98" />
                    <SPLIT distance="550" swimtime="00:06:14.69" />
                    <SPLIT distance="600" swimtime="00:06:49.54" />
                    <SPLIT distance="650" swimtime="00:07:25.24" />
                    <SPLIT distance="700" swimtime="00:08:00.31" />
                    <SPLIT distance="750" swimtime="00:08:34.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="445" swimtime="00:02:26.59" resultid="8907" heatid="10479" lane="3" entrytime="00:02:25.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.69" />
                    <SPLIT distance="100" swimtime="00:01:12.08" />
                    <SPLIT distance="150" swimtime="00:01:49.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="522" swimtime="00:05:01.01" resultid="8908" heatid="10523" lane="1" entrytime="00:05:04.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                    <SPLIT distance="100" swimtime="00:01:08.68" />
                    <SPLIT distance="150" swimtime="00:01:48.27" />
                    <SPLIT distance="200" swimtime="00:02:26.43" />
                    <SPLIT distance="250" swimtime="00:03:11.34" />
                    <SPLIT distance="300" swimtime="00:03:55.08" />
                    <SPLIT distance="350" swimtime="00:04:29.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1257" points="582" swimtime="00:17:22.80" resultid="8909" heatid="10635" lane="6" entrytime="00:17:25.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.82" />
                    <SPLIT distance="100" swimtime="00:01:03.31" />
                    <SPLIT distance="150" swimtime="00:01:36.94" />
                    <SPLIT distance="200" swimtime="00:02:11.27" />
                    <SPLIT distance="250" swimtime="00:02:46.04" />
                    <SPLIT distance="300" swimtime="00:03:21.28" />
                    <SPLIT distance="350" swimtime="00:03:56.20" />
                    <SPLIT distance="400" swimtime="00:04:31.22" />
                    <SPLIT distance="450" swimtime="00:05:06.48" />
                    <SPLIT distance="500" swimtime="00:05:41.25" />
                    <SPLIT distance="550" swimtime="00:06:16.82" />
                    <SPLIT distance="600" swimtime="00:06:51.89" />
                    <SPLIT distance="650" swimtime="00:07:27.50" />
                    <SPLIT distance="700" swimtime="00:08:02.75" />
                    <SPLIT distance="750" swimtime="00:08:38.27" />
                    <SPLIT distance="800" swimtime="00:09:13.64" />
                    <SPLIT distance="850" swimtime="00:09:48.52" />
                    <SPLIT distance="900" swimtime="00:10:23.33" />
                    <SPLIT distance="950" swimtime="00:10:59.21" />
                    <SPLIT distance="1000" swimtime="00:11:34.38" />
                    <SPLIT distance="1050" swimtime="00:12:10.29" />
                    <SPLIT distance="1100" swimtime="00:12:45.60" />
                    <SPLIT distance="1150" swimtime="00:13:21.20" />
                    <SPLIT distance="1200" swimtime="00:13:56.48" />
                    <SPLIT distance="1250" swimtime="00:14:29.46" />
                    <SPLIT distance="1300" swimtime="00:15:04.92" />
                    <SPLIT distance="1350" swimtime="00:15:40.62" />
                    <SPLIT distance="1400" swimtime="00:16:15.85" />
                    <SPLIT distance="1450" swimtime="00:16:50.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="477" swimtime="00:02:25.85" resultid="8910" heatid="10651" lane="6" entrytime="00:02:24.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                    <SPLIT distance="100" swimtime="00:01:10.78" />
                    <SPLIT distance="150" swimtime="00:01:54.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1357" points="567" swimtime="00:04:25.88" resultid="8911" heatid="10723" lane="4" entrytime="00:04:27.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                    <SPLIT distance="100" swimtime="00:01:03.24" />
                    <SPLIT distance="150" swimtime="00:01:37.60" />
                    <SPLIT distance="200" swimtime="00:02:12.23" />
                    <SPLIT distance="250" swimtime="00:02:46.44" />
                    <SPLIT distance="300" swimtime="00:03:19.92" />
                    <SPLIT distance="350" swimtime="00:03:54.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Cecilia Zampieri" birthdate="2010-09-17" gender="F" nation="BRA" license="421899" swrid="5820335" athleteid="9058" externalid="421899">
              <RESULTS>
                <RESULT comment="SW 6.4 - A virada não foi iniciada após a conclusão do movimento de braço, após sair da posição de costas.  (Horário: 9:00), Na volta dos 100m." eventid="1063" status="DSQ" swimtime="00:03:09.24" resultid="9059" heatid="10469" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="285" swimtime="00:01:18.55" resultid="9060" heatid="10524" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="248" swimtime="00:00:42.70" resultid="9061" heatid="10676" lane="5" />
                <RESULT eventid="1365" points="231" swimtime="00:01:33.07" resultid="9062" heatid="10728" lane="0" entrytime="00:01:29.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Kozera Chiarato" birthdate="2010-05-28" gender="M" nation="BRA" license="406722" swrid="5717275" athleteid="9010" externalid="406722">
              <RESULTS>
                <RESULT eventid="1123" points="323" swimtime="00:10:58.62" resultid="9011" heatid="10516" lane="2" entrytime="00:11:02.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.42" />
                    <SPLIT distance="100" swimtime="00:01:12.69" />
                    <SPLIT distance="150" swimtime="00:01:53.23" />
                    <SPLIT distance="200" swimtime="00:02:35.29" />
                    <SPLIT distance="250" swimtime="00:03:17.66" />
                    <SPLIT distance="300" swimtime="00:04:00.99" />
                    <SPLIT distance="350" swimtime="00:04:43.85" />
                    <SPLIT distance="400" swimtime="00:05:26.31" />
                    <SPLIT distance="450" swimtime="00:06:09.06" />
                    <SPLIT distance="500" swimtime="00:06:51.50" />
                    <SPLIT distance="550" swimtime="00:07:33.55" />
                    <SPLIT distance="600" swimtime="00:08:15.60" />
                    <SPLIT distance="650" swimtime="00:08:57.77" />
                    <SPLIT distance="700" swimtime="00:09:39.68" />
                    <SPLIT distance="750" swimtime="00:10:20.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="356" swimtime="00:00:31.41" resultid="9012" heatid="10504" lane="5" entrytime="00:00:33.21" entrycourse="LCM" />
                <RESULT eventid="1171" points="254" swimtime="00:02:54.11" resultid="9013" heatid="10556" lane="8" entrytime="00:03:03.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                    <SPLIT distance="100" swimtime="00:01:15.37" />
                    <SPLIT distance="150" swimtime="00:02:02.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="342" swimtime="00:01:06.29" resultid="9014" heatid="10545" lane="7" entrytime="00:01:04.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="287" swimtime="00:02:52.80" resultid="9015" heatid="10648" lane="8" entrytime="00:02:53.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                    <SPLIT distance="100" swimtime="00:01:24.75" />
                    <SPLIT distance="150" swimtime="00:02:16.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1341" points="328" swimtime="00:01:11.64" resultid="9016" heatid="10707" lane="7" entrytime="00:01:13.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Vitor Navarro Zanini" birthdate="2008-06-30" gender="M" nation="BRA" license="369415" swrid="5600273" athleteid="8958" externalid="369415">
              <RESULTS>
                <RESULT eventid="1087" points="364" swimtime="00:02:55.70" resultid="8959" heatid="10490" lane="6" entrytime="00:02:55.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                    <SPLIT distance="100" swimtime="00:01:20.75" />
                    <SPLIT distance="150" swimtime="00:02:06.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="432" swimtime="00:00:34.32" resultid="8960" heatid="10573" lane="4" entrytime="00:00:35.54" entrycourse="LCM" />
                <RESULT eventid="1219" points="400" swimtime="00:01:17.16" resultid="8961" heatid="10596" lane="6" entrytime="00:01:18.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="389" swimtime="00:02:19.68" resultid="8962" heatid="10669" lane="4" entrytime="00:02:18.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="100" swimtime="00:01:07.74" />
                    <SPLIT distance="150" swimtime="00:01:44.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaylane" lastname="Marques Ferreira" birthdate="2010-03-06" gender="F" nation="BRA" license="391146" swrid="5600211" athleteid="8984" externalid="391146">
              <RESULTS>
                <RESULT eventid="1095" points="397" swimtime="00:00:33.23" resultid="8985" heatid="10497" lane="7" entrytime="00:00:34.60" entrycourse="LCM" />
                <RESULT eventid="1163" points="247" swimtime="00:03:13.96" resultid="8986" heatid="10554" lane="9" entrytime="00:03:19.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                    <SPLIT distance="100" swimtime="00:01:25.95" />
                    <SPLIT distance="150" swimtime="00:02:26.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="258" swimtime="00:03:17.96" resultid="8987" heatid="10640" lane="9" entrytime="00:03:28.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                    <SPLIT distance="100" swimtime="00:01:25.47" />
                    <SPLIT distance="150" swimtime="00:02:34.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="269" swimtime="00:02:53.83" resultid="8988" heatid="10655" lane="9" entrytime="00:02:45.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                    <SPLIT distance="100" swimtime="00:01:21.67" />
                    <SPLIT distance="150" swimtime="00:02:10.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="251" swimtime="00:06:12.77" resultid="8989" heatid="10712" lane="3" entrytime="00:06:22.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.88" />
                    <SPLIT distance="100" swimtime="00:01:25.91" />
                    <SPLIT distance="150" swimtime="00:02:15.47" />
                    <SPLIT distance="200" swimtime="00:03:05.43" />
                    <SPLIT distance="250" swimtime="00:03:55.08" />
                    <SPLIT distance="300" swimtime="00:04:46.15" />
                    <SPLIT distance="350" swimtime="00:05:29.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="344" swimtime="00:01:18.68" resultid="8990" heatid="10701" lane="7" entrytime="00:01:20.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monike" lastname="Lemos Carvalho" birthdate="2008-03-28" gender="F" nation="BRA" license="307796" swrid="5600199" athleteid="8963" externalid="307796">
              <RESULTS>
                <RESULT eventid="1115" points="388" swimtime="00:21:02.00" resultid="8964" heatid="10512" lane="2" entrytime="00:21:03.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                    <SPLIT distance="100" swimtime="00:01:14.13" />
                    <SPLIT distance="150" swimtime="00:01:51.75" />
                    <SPLIT distance="200" swimtime="00:02:30.41" />
                    <SPLIT distance="250" swimtime="00:03:10.38" />
                    <SPLIT distance="300" swimtime="00:03:51.67" />
                    <SPLIT distance="350" swimtime="00:04:33.36" />
                    <SPLIT distance="400" swimtime="00:05:16.44" />
                    <SPLIT distance="450" swimtime="00:05:59.26" />
                    <SPLIT distance="500" swimtime="00:06:42.49" />
                    <SPLIT distance="550" swimtime="00:07:25.60" />
                    <SPLIT distance="600" swimtime="00:08:09.09" />
                    <SPLIT distance="650" swimtime="00:08:52.20" />
                    <SPLIT distance="700" swimtime="00:09:34.88" />
                    <SPLIT distance="750" swimtime="00:10:17.76" />
                    <SPLIT distance="800" swimtime="00:11:00.26" />
                    <SPLIT distance="850" swimtime="00:11:43.38" />
                    <SPLIT distance="900" swimtime="00:12:26.74" />
                    <SPLIT distance="950" swimtime="00:13:10.18" />
                    <SPLIT distance="1000" swimtime="00:13:53.76" />
                    <SPLIT distance="1050" swimtime="00:14:37.19" />
                    <SPLIT distance="1100" swimtime="00:15:21.19" />
                    <SPLIT distance="1150" swimtime="00:16:04.49" />
                    <SPLIT distance="1200" swimtime="00:16:48.02" />
                    <SPLIT distance="1250" swimtime="00:17:31.14" />
                    <SPLIT distance="1300" swimtime="00:18:13.95" />
                    <SPLIT distance="1350" swimtime="00:18:57.17" />
                    <SPLIT distance="1400" swimtime="00:19:39.49" />
                    <SPLIT distance="1450" swimtime="00:20:21.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="347" swimtime="00:02:55.22" resultid="8965" heatid="10470" lane="5" entrytime="00:02:57.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="428" swimtime="00:10:43.11" resultid="8966" heatid="10633" lane="5" entrytime="00:11:01.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                    <SPLIT distance="100" swimtime="00:01:11.58" />
                    <SPLIT distance="150" swimtime="00:01:49.82" />
                    <SPLIT distance="200" swimtime="00:02:28.65" />
                    <SPLIT distance="250" swimtime="00:03:08.59" />
                    <SPLIT distance="300" swimtime="00:03:49.63" />
                    <SPLIT distance="350" swimtime="00:04:30.31" />
                    <SPLIT distance="400" swimtime="00:05:11.25" />
                    <SPLIT distance="450" swimtime="00:05:52.91" />
                    <SPLIT distance="500" swimtime="00:06:34.69" />
                    <SPLIT distance="550" swimtime="00:07:16.31" />
                    <SPLIT distance="600" swimtime="00:07:59.04" />
                    <SPLIT distance="650" swimtime="00:08:40.92" />
                    <SPLIT distance="700" swimtime="00:09:22.39" />
                    <SPLIT distance="750" swimtime="00:10:03.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="505" swimtime="00:02:20.92" resultid="8967" heatid="10659" lane="3" entrytime="00:02:21.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                    <SPLIT distance="100" swimtime="00:01:07.65" />
                    <SPLIT distance="150" swimtime="00:01:44.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="422" swimtime="00:05:13.60" resultid="8968" heatid="10714" lane="4" entrytime="00:05:12.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                    <SPLIT distance="100" swimtime="00:01:11.57" />
                    <SPLIT distance="150" swimtime="00:01:50.48" />
                    <SPLIT distance="200" swimtime="00:02:31.00" />
                    <SPLIT distance="250" swimtime="00:03:12.06" />
                    <SPLIT distance="300" swimtime="00:03:53.07" />
                    <SPLIT distance="350" swimtime="00:04:33.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="377" swimtime="00:01:19.04" resultid="8969" heatid="10731" lane="1" entrytime="00:01:16.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduarda" lastname="Azevedo Birsneek" birthdate="2010-03-31" gender="F" nation="BRA" license="391145" swrid="5389427" athleteid="8977" externalid="391145">
              <RESULTS>
                <RESULT eventid="1095" points="166" swimtime="00:00:44.38" resultid="8978" heatid="10495" lane="7" entrytime="00:00:47.45" entrycourse="LCM" />
                <RESULT eventid="1063" points="203" swimtime="00:03:29.21" resultid="8979" heatid="10470" lane="0" entrytime="00:03:15.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="220" swimtime="00:00:44.49" resultid="8980" heatid="10678" lane="8" entrytime="00:00:43.93" entrycourse="LCM" />
                <RESULT eventid="1265" points="192" swimtime="00:03:38.37" resultid="8981" heatid="10639" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.66" />
                    <SPLIT distance="100" swimtime="00:01:38.84" />
                    <SPLIT distance="150" swimtime="00:02:48.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1333" points="136" swimtime="00:01:47.09" resultid="8982" heatid="10699" lane="5" entrytime="00:01:45.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="220" swimtime="00:01:34.60" resultid="8983" heatid="10727" lane="7" entrytime="00:01:34.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Rodrigues Galvao" birthdate="2007-04-19" gender="M" nation="BRA" license="376586" swrid="5600247" athleteid="8890" externalid="376586">
              <RESULTS>
                <RESULT eventid="1103" points="509" swimtime="00:00:27.89" resultid="8891" heatid="10508" lane="9" entrytime="00:00:27.64" entrycourse="LCM" />
                <RESULT eventid="1171" points="372" swimtime="00:02:33.31" resultid="8892" heatid="10557" lane="6" entrytime="00:02:33.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.19" />
                    <SPLIT distance="100" swimtime="00:01:10.12" />
                    <SPLIT distance="150" swimtime="00:01:51.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="489" swimtime="00:00:26.53" resultid="8893" heatid="10626" lane="7" entrytime="00:00:25.92" entrycourse="LCM" />
                <RESULT eventid="1341" points="502" swimtime="00:01:02.18" resultid="8894" heatid="10710" lane="1" entrytime="00:01:03.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Luiza Rimbano De Jesus" birthdate="2008-09-02" gender="F" nation="BRA" license="366819" swrid="5653297" athleteid="8996" externalid="366819">
              <RESULTS>
                <RESULT eventid="1179" points="426" swimtime="00:00:38.73" resultid="8997" heatid="10564" lane="3" entrytime="00:00:37.45" entrycourse="LCM" />
                <RESULT eventid="1147" points="556" swimtime="00:01:02.88" resultid="8998" heatid="10534" lane="6" entrytime="00:01:02.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="552" swimtime="00:00:28.77" resultid="8999" heatid="10609" lane="3" entrytime="00:00:28.16" entrycourse="LCM" />
                <RESULT eventid="1211" points="351" swimtime="00:01:30.88" resultid="9000" heatid="10587" lane="7" entrytime="00:01:25.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1281" points="447" swimtime="00:02:26.75" resultid="9001" heatid="10659" lane="9" entrytime="00:02:23.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                    <SPLIT distance="100" swimtime="00:01:08.95" />
                    <SPLIT distance="150" swimtime="00:01:47.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1365" points="357" swimtime="00:01:20.53" resultid="9002" heatid="10729" lane="5" entrytime="00:01:21.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lauren" lastname="Dziura" birthdate="2010-01-11" gender="F" nation="BRA" license="369416" swrid="5588668" athleteid="8926" externalid="369416">
              <RESULTS>
                <RESULT eventid="1115" points="432" swimtime="00:20:16.88" resultid="8927" heatid="10512" lane="5" entrytime="00:20:28.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                    <SPLIT distance="100" swimtime="00:01:15.48" />
                    <SPLIT distance="150" swimtime="00:01:55.29" />
                    <SPLIT distance="200" swimtime="00:02:35.27" />
                    <SPLIT distance="250" swimtime="00:03:15.11" />
                    <SPLIT distance="300" swimtime="00:03:55.54" />
                    <SPLIT distance="350" swimtime="00:04:35.70" />
                    <SPLIT distance="400" swimtime="00:05:15.98" />
                    <SPLIT distance="450" swimtime="00:05:56.21" />
                    <SPLIT distance="500" swimtime="00:06:36.72" />
                    <SPLIT distance="550" swimtime="00:07:16.62" />
                    <SPLIT distance="600" swimtime="00:07:57.10" />
                    <SPLIT distance="650" swimtime="00:08:38.18" />
                    <SPLIT distance="700" swimtime="00:09:18.62" />
                    <SPLIT distance="750" swimtime="00:09:59.65" />
                    <SPLIT distance="800" swimtime="00:10:41.48" />
                    <SPLIT distance="850" swimtime="00:11:22.94" />
                    <SPLIT distance="900" swimtime="00:12:03.70" />
                    <SPLIT distance="950" swimtime="00:12:44.74" />
                    <SPLIT distance="1000" swimtime="00:13:25.48" />
                    <SPLIT distance="1050" swimtime="00:14:06.29" />
                    <SPLIT distance="1100" swimtime="00:14:48.16" />
                    <SPLIT distance="1150" swimtime="00:15:29.10" />
                    <SPLIT distance="1200" swimtime="00:16:11.02" />
                    <SPLIT distance="1250" swimtime="00:16:51.72" />
                    <SPLIT distance="1300" swimtime="00:17:33.80" />
                    <SPLIT distance="1350" swimtime="00:18:15.83" />
                    <SPLIT distance="1400" swimtime="00:18:57.90" />
                    <SPLIT distance="1450" swimtime="00:19:38.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="323" swimtime="00:06:25.02" resultid="8928" heatid="10519" lane="8" entrytime="00:06:18.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.35" />
                    <SPLIT distance="100" swimtime="00:01:33.92" />
                    <SPLIT distance="150" swimtime="00:02:24.39" />
                    <SPLIT distance="200" swimtime="00:03:13.47" />
                    <SPLIT distance="250" swimtime="00:04:10.38" />
                    <SPLIT distance="300" swimtime="00:05:04.52" />
                    <SPLIT distance="350" swimtime="00:05:45.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="423" swimtime="00:10:45.81" resultid="8929" heatid="10632" lane="9" entrytime="00:10:54.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.95" />
                    <SPLIT distance="100" swimtime="00:01:13.63" />
                    <SPLIT distance="150" swimtime="00:01:53.67" />
                    <SPLIT distance="200" swimtime="00:02:34.73" />
                    <SPLIT distance="250" swimtime="00:03:15.18" />
                    <SPLIT distance="300" swimtime="00:03:56.44" />
                    <SPLIT distance="350" swimtime="00:04:37.28" />
                    <SPLIT distance="400" swimtime="00:05:19.04" />
                    <SPLIT distance="450" swimtime="00:06:00.95" />
                    <SPLIT distance="500" swimtime="00:06:42.31" />
                    <SPLIT distance="550" swimtime="00:07:23.34" />
                    <SPLIT distance="600" swimtime="00:08:04.73" />
                    <SPLIT distance="650" swimtime="00:08:45.72" />
                    <SPLIT distance="700" swimtime="00:09:27.35" />
                    <SPLIT distance="750" swimtime="00:10:06.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="289" swimtime="00:00:40.62" resultid="8930" heatid="10675" lane="5" />
                <RESULT eventid="1265" points="332" swimtime="00:03:01.96" resultid="8931" heatid="10641" lane="2" entrytime="00:02:59.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.58" />
                    <SPLIT distance="100" swimtime="00:01:30.32" />
                    <SPLIT distance="150" swimtime="00:02:24.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1349" points="416" swimtime="00:05:15.29" resultid="8932" heatid="10715" lane="0" entrytime="00:05:11.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.81" />
                    <SPLIT distance="100" swimtime="00:01:14.23" />
                    <SPLIT distance="150" swimtime="00:01:54.31" />
                    <SPLIT distance="200" swimtime="00:02:34.01" />
                    <SPLIT distance="250" swimtime="00:03:15.45" />
                    <SPLIT distance="300" swimtime="00:03:56.08" />
                    <SPLIT distance="350" swimtime="00:04:36.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stella" lastname="Magalhaes Birnbaum" birthdate="2009-05-14" gender="F" nation="BRA" license="399684" swrid="5653298" athleteid="9063" externalid="399684">
              <RESULTS>
                <RESULT eventid="1095" points="228" swimtime="00:00:39.95" resultid="9064" heatid="10496" lane="1" entrytime="00:00:39.45" entrycourse="LCM" />
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 19:12)" eventid="1179" status="DSQ" swimtime="00:00:50.75" resultid="9065" heatid="10561" lane="1" />
                <RESULT eventid="1227" points="318" swimtime="00:00:34.56" resultid="9066" heatid="10604" lane="4" entrytime="00:00:31.72" entrycourse="LCM" />
                <RESULT eventid="1297" points="357" swimtime="00:00:37.83" resultid="9067" heatid="10679" lane="1" entrytime="00:00:38.87" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Lemes Luis" birthdate="2011-11-10" gender="M" nation="BRA" license="421440" swrid="5810967" athleteid="9038" externalid="421440">
              <RESULTS>
                <RESULT eventid="1123" points="313" swimtime="00:11:05.34" resultid="9039" heatid="10516" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.64" />
                    <SPLIT distance="100" swimtime="00:01:17.71" />
                    <SPLIT distance="150" swimtime="00:01:59.89" />
                    <SPLIT distance="200" swimtime="00:02:42.93" />
                    <SPLIT distance="250" swimtime="00:03:25.34" />
                    <SPLIT distance="300" swimtime="00:04:07.56" />
                    <SPLIT distance="350" swimtime="00:04:50.39" />
                    <SPLIT distance="400" swimtime="00:05:33.27" />
                    <SPLIT distance="450" swimtime="00:06:15.66" />
                    <SPLIT distance="500" swimtime="00:06:57.67" />
                    <SPLIT distance="550" swimtime="00:07:39.52" />
                    <SPLIT distance="600" swimtime="00:08:21.67" />
                    <SPLIT distance="650" swimtime="00:09:03.61" />
                    <SPLIT distance="700" swimtime="00:09:45.87" />
                    <SPLIT distance="750" swimtime="00:10:25.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="166" swimtime="00:00:40.50" resultid="9040" heatid="10500" lane="5" />
                <RESULT eventid="1155" points="280" swimtime="00:01:10.88" resultid="9041" heatid="10541" lane="8" entrytime="00:01:11.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="255" swimtime="00:00:32.97" resultid="9042" heatid="10612" lane="0" />
                <RESULT eventid="1219" points="189" swimtime="00:01:39.06" resultid="9043" heatid="10591" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1331" points="424" swimtime="00:04:35.14" resultid="9077" heatid="10698" lane="2" entrytime="00:04:34.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                    <SPLIT distance="100" swimtime="00:01:09.74" />
                    <SPLIT distance="150" swimtime="00:01:47.32" />
                    <SPLIT distance="200" swimtime="00:02:29.39" />
                    <SPLIT distance="250" swimtime="00:02:59.35" />
                    <SPLIT distance="300" swimtime="00:03:32.96" />
                    <SPLIT distance="350" swimtime="00:04:02.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8919" number="1" />
                    <RELAYPOSITION athleteid="8958" number="2" />
                    <RELAYPOSITION athleteid="8890" number="3" />
                    <RELAYPOSITION athleteid="8940" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1399" points="464" swimtime="00:04:03.11" resultid="9079" heatid="10753" lane="6" entrytime="00:03:51.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.89" />
                    <SPLIT distance="100" swimtime="00:00:58.89" />
                    <SPLIT distance="150" swimtime="00:01:28.73" />
                    <SPLIT distance="200" swimtime="00:02:01.88" />
                    <SPLIT distance="250" swimtime="00:02:33.17" />
                    <SPLIT distance="300" swimtime="00:03:06.15" />
                    <SPLIT distance="350" swimtime="00:03:33.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8890" number="1" />
                    <RELAYPOSITION athleteid="8940" number="2" />
                    <RELAYPOSITION athleteid="8958" number="3" />
                    <RELAYPOSITION athleteid="8919" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1325" points="285" swimtime="00:05:13.95" resultid="9078" heatid="10695" lane="7" entrytime="00:05:04.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                    <SPLIT distance="100" swimtime="00:01:15.13" />
                    <SPLIT distance="150" swimtime="00:01:52.70" />
                    <SPLIT distance="200" swimtime="00:02:35.55" />
                    <SPLIT distance="250" swimtime="00:03:16.62" />
                    <SPLIT distance="300" swimtime="00:04:04.87" />
                    <SPLIT distance="350" swimtime="00:04:37.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8970" number="1" />
                    <RELAYPOSITION athleteid="9003" number="2" />
                    <RELAYPOSITION athleteid="8991" number="3" />
                    <RELAYPOSITION athleteid="9038" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1395" points="366" swimtime="00:04:23.05" resultid="9080" heatid="10751" lane="6" entrytime="00:04:23.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.37" />
                    <SPLIT distance="100" swimtime="00:01:02.94" />
                    <SPLIT distance="150" swimtime="00:01:32.21" />
                    <SPLIT distance="200" swimtime="00:02:04.39" />
                    <SPLIT distance="250" swimtime="00:02:36.00" />
                    <SPLIT distance="300" swimtime="00:03:10.44" />
                    <SPLIT distance="350" swimtime="00:03:43.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8945" number="1" />
                    <RELAYPOSITION athleteid="8933" number="2" />
                    <RELAYPOSITION athleteid="9010" number="3" />
                    <RELAYPOSITION athleteid="9024" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="F" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1321" points="379" swimtime="00:05:17.17" resultid="9073" heatid="10692" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.77" />
                    <SPLIT distance="100" swimtime="00:01:18.79" />
                    <SPLIT distance="150" swimtime="00:01:59.35" />
                    <SPLIT distance="200" swimtime="00:02:48.73" />
                    <SPLIT distance="250" swimtime="00:03:25.65" />
                    <SPLIT distance="300" swimtime="00:04:14.22" />
                    <SPLIT distance="350" swimtime="00:04:43.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8963" number="1" />
                    <RELAYPOSITION athleteid="8895" number="2" />
                    <RELAYPOSITION athleteid="8898" number="3" />
                    <RELAYPOSITION athleteid="8996" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="F" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1317" points="339" swimtime="00:05:29.20" resultid="9074" heatid="10690" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                    <SPLIT distance="100" swimtime="00:01:26.38" />
                    <SPLIT distance="150" swimtime="00:02:02.87" />
                    <SPLIT distance="200" swimtime="00:02:46.35" />
                    <SPLIT distance="250" swimtime="00:03:22.02" />
                    <SPLIT distance="300" swimtime="00:04:09.35" />
                    <SPLIT distance="350" swimtime="00:04:46.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8926" number="1" />
                    <RELAYPOSITION athleteid="8870" number="2" />
                    <RELAYPOSITION athleteid="8984" number="3" />
                    <RELAYPOSITION athleteid="9058" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1385" points="334" swimtime="00:04:59.56" resultid="9075" heatid="10745" lane="0">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                    <SPLIT distance="100" swimtime="00:01:09.92" />
                    <SPLIT distance="150" swimtime="00:01:48.72" />
                    <SPLIT distance="200" swimtime="00:02:31.48" />
                    <SPLIT distance="250" swimtime="00:03:06.93" />
                    <SPLIT distance="300" swimtime="00:03:49.60" />
                    <SPLIT distance="350" swimtime="00:04:22.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="8870" number="1" />
                    <RELAYPOSITION athleteid="9058" number="2" />
                    <RELAYPOSITION athleteid="8984" number="3" />
                    <RELAYPOSITION athleteid="8926" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1383" points="307" swimtime="00:05:07.99" resultid="9076" heatid="10744" lane="1" entrytime="00:05:10.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                    <SPLIT distance="100" swimtime="00:01:15.16" />
                    <SPLIT distance="150" swimtime="00:01:53.44" />
                    <SPLIT distance="200" swimtime="00:02:37.41" />
                    <SPLIT distance="250" swimtime="00:03:12.45" />
                    <SPLIT distance="300" swimtime="00:03:52.16" />
                    <SPLIT distance="350" swimtime="00:04:27.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="9044" number="1" />
                    <RELAYPOSITION athleteid="9031" number="2" />
                    <RELAYPOSITION athleteid="9017" number="3" />
                    <RELAYPOSITION athleteid="8883" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
