<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.77033">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Campo Mourão" name="Torneio Regional da 2ª Região (Pré-Mirim/Sênior)" course="SCM" deadline="2023-03-14" entrystartdate="2023-03-07" entrytype="INVITATION" hostclub="Fundação de Esportes de Campo Mourão" hostclub.url="https://campomourao.atende.net/subportal/fundacao-de-esportes" number="37074" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/evento/natacao/37074" startmethod="2" timing="AUTOMATIC" withdrawuntil="2023-03-15" state="PR" nation="BRA" maxentriesathlete="6">
      <AGEDATE value="2023-01-01" type="YEAR" />
      <POOL name="Complexo Esportivo Roberto Brzezinski" lanemin="2" lanemax="7" />
      <FACILITY city="Campo Mourão" name="Complexo Esportivo Roberto Brzezinski" nation="BRA" state="PR" street="Rua Miguel Luís Pereira" street2="Bela Vista" zip="87302-140" />
      <POINTTABLE pointtableid="3015" name="FINA Point Scoring" version="2022" />
      <QUALIFY from="2022-03-18" until="2022-03-18" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99252-0598" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99252-0598" street="Avenida do Batel, 1230" street2="Sala 202" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2023-03-18" daytime="09:10" number="1" teamleadermeeting="09:00" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="1061" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1062" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5394" />
                    <RANKING order="2" place="2" resultid="5410" />
                    <RANKING order="3" place="3" resultid="5421" />
                    <RANKING order="4" place="4" resultid="5407" />
                    <RANKING order="5" place="5" resultid="5164" />
                    <RANKING order="6" place="6" resultid="5364" />
                    <RANKING order="7" place="7" resultid="5430" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1063" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5131" />
                    <RANKING order="2" place="2" resultid="5146" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4850" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4851" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1064" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1065" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5399" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5126" />
                    <RANKING order="2" place="2" resultid="5437" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4852" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1067" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1068" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5241" />
                    <RANKING order="2" place="2" resultid="5343" />
                    <RANKING order="3" place="3" resultid="5236" />
                    <RANKING order="4" place="4" resultid="5002" />
                    <RANKING order="5" place="-1" resultid="4984" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1070" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5015" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1072" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1073" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1074" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4853" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1075" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1076" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5108" />
                    <RANKING order="2" place="2" resultid="5382" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1077" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5102" />
                    <RANKING order="2" place="2" resultid="5157" />
                    <RANKING order="3" place="-1" resultid="5417" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1078" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5046" />
                    <RANKING order="2" place="2" resultid="4996" />
                    <RANKING order="3" place="3" resultid="5067" />
                    <RANKING order="4" place="4" resultid="5291" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1079" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4978" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1080" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5070" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1081" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5056" />
                    <RANKING order="2" place="2" resultid="5355" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5491" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4854" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4855" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4856" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1085" gender="M" number="6" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1086" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5469" />
                    <RANKING order="2" place="2" resultid="5288" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4857" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1087" gender="F" number="7" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1088" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5227" />
                    <RANKING order="2" place="2" resultid="5458" />
                    <RANKING order="3" place="3" resultid="5465" />
                    <RANKING order="4" place="-1" resultid="5530" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1089" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5168" />
                    <RANKING order="2" place="2" resultid="5425" />
                    <RANKING order="3" place="3" resultid="5141" />
                    <RANKING order="4" place="4" resultid="5335" />
                    <RANKING order="5" place="5" resultid="5433" />
                    <RANKING order="6" place="6" resultid="5374" />
                    <RANKING order="7" place="7" resultid="5211" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4858" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4859" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1090" gender="M" number="8" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1091" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5262" />
                    <RANKING order="2" place="2" resultid="5528" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1092" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5179" />
                    <RANKING order="2" place="2" resultid="5309" />
                    <RANKING order="3" place="3" resultid="5445" />
                    <RANKING order="4" place="4" resultid="5467" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4860" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1093" gender="F" number="9" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1094" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5163" />
                    <RANKING order="2" place="2" resultid="5363" />
                    <RANKING order="3" place="3" resultid="5429" />
                    <RANKING order="4" place="4" resultid="5216" />
                    <RANKING order="5" place="5" resultid="5406" />
                    <RANKING order="6" place="6" resultid="5522" />
                    <RANKING order="7" place="7" resultid="5455" />
                    <RANKING order="8" place="8" resultid="5251" />
                    <RANKING order="9" place="-1" resultid="5267" />
                    <RANKING order="10" place="-1" resultid="5526" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1095" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5275" />
                    <RANKING order="2" place="2" resultid="5283" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4861" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4862" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1096" gender="M" number="10" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1097" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5190" />
                    <RANKING order="2" place="2" resultid="5173" />
                    <RANKING order="3" place="3" resultid="5398" />
                    <RANKING order="4" place="4" resultid="5537" />
                    <RANKING order="5" place="5" resultid="5184" />
                    <RANKING order="6" place="6" resultid="5196" />
                    <RANKING order="7" place="7" resultid="5386" />
                    <RANKING order="8" place="8" resultid="5524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5390" />
                    <RANKING order="2" place="2" resultid="5414" />
                    <RANKING order="3" place="3" resultid="5476" />
                    <RANKING order="4" place="4" resultid="5271" />
                    <RANKING order="5" place="5" resultid="5532" />
                    <RANKING order="6" place="-1" resultid="5487" />
                    <RANKING order="7" place="-1" resultid="5122" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4863" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4864" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4865" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1099" gender="F" number="11" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1100" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1101" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5082" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1103" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5331" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1104" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5494" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1105" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1106" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4866" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1107" gender="M" number="12" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1108" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1109" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5418" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1110" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5097" />
                    <RANKING order="2" place="2" resultid="5351" />
                    <RANKING order="3" place="3" resultid="5347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1111" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5511" />
                    <RANKING order="2" place="2" resultid="5232" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1112" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5060" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1113" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1114" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5339" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4867" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4868" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1115" gender="F" number="13" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1116" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5402" />
                    <RANKING order="2" place="2" resultid="5371" />
                    <RANKING order="3" place="3" resultid="5441" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1117" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5021" />
                    <RANKING order="2" place="2" resultid="5426" />
                    <RANKING order="3" place="3" resultid="5142" />
                    <RANKING order="4" place="4" resultid="5336" />
                    <RANKING order="5" place="5" resultid="5434" />
                    <RANKING order="6" place="6" resultid="5480" />
                    <RANKING order="7" place="7" resultid="5461" />
                    <RANKING order="8" place="8" resultid="5212" />
                    <RANKING order="9" place="9" resultid="5359" />
                    <RANKING order="10" place="10" resultid="5375" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4869" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4870" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4871" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1118" gender="M" number="14" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1119" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5255" />
                    <RANKING order="2" place="2" resultid="5300" />
                    <RANKING order="3" place="3" resultid="5263" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1120" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5180" />
                    <RANKING order="2" place="2" resultid="5222" />
                    <RANKING order="3" place="3" resultid="5317" />
                    <RANKING order="4" place="4" resultid="5279" />
                    <RANKING order="5" place="5" resultid="5310" />
                    <RANKING order="6" place="6" resultid="5304" />
                    <RANKING order="7" place="7" resultid="5446" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4872" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4873" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1121" gender="F" number="15" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1122" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5206" />
                    <RANKING order="2" place="2" resultid="5217" />
                    <RANKING order="3" place="3" resultid="5367" />
                    <RANKING order="4" place="4" resultid="5252" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1123" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5132" />
                    <RANKING order="2" place="2" resultid="5147" />
                    <RANKING order="3" place="3" resultid="5276" />
                    <RANKING order="4" place="4" resultid="5323" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4874" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4875" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1124" gender="M" number="16" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1125" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5191" />
                    <RANKING order="2" place="2" resultid="5174" />
                    <RANKING order="3" place="3" resultid="5152" />
                    <RANKING order="4" place="4" resultid="5387" />
                    <RANKING order="5" place="5" resultid="5197" />
                    <RANKING order="6" place="6" resultid="5448" />
                    <RANKING order="7" place="7" resultid="5185" />
                    <RANKING order="8" place="8" resultid="5313" />
                    <RANKING order="9" place="9" resultid="5538" />
                    <RANKING order="10" place="10" resultid="5137" />
                    <RANKING order="11" place="11" resultid="5378" />
                    <RANKING order="12" place="12" resultid="5296" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5415" />
                    <RANKING order="2" place="2" resultid="5201" />
                    <RANKING order="3" place="3" resultid="5391" />
                    <RANKING order="4" place="4" resultid="5438" />
                    <RANKING order="5" place="5" resultid="5008" />
                    <RANKING order="6" place="6" resultid="5477" />
                    <RANKING order="7" place="7" resultid="5272" />
                    <RANKING order="8" place="8" resultid="5473" />
                    <RANKING order="9" place="9" resultid="5483" />
                    <RANKING order="10" place="-1" resultid="5123" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4876" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4877" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4878" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4879" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1127" gender="F" number="17" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1128" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5242" />
                    <RANKING order="2" place="2" resultid="4985" />
                    <RANKING order="3" place="3" resultid="5003" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1129" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5087" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1130" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5092" />
                    <RANKING order="2" place="2" resultid="5062" />
                    <RANKING order="3" place="3" resultid="5016" />
                    <RANKING order="4" place="4" resultid="5247" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1131" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4990" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1132" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1133" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5058" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1134" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5052" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4880" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4881" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1135" gender="M" number="18" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1136" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5118" />
                    <RANKING order="2" place="2" resultid="5327" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1137" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5076" />
                    <RANKING order="2" place="2" resultid="5103" />
                    <RANKING order="3" place="3" resultid="5513" />
                    <RANKING order="4" place="4" resultid="5158" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1138" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5031" />
                    <RANKING order="2" place="2" resultid="5036" />
                    <RANKING order="3" place="3" resultid="4997" />
                    <RANKING order="4" place="4" resultid="5285" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1139" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5233" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1140" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5026" />
                    <RANKING order="2" place="2" resultid="5061" />
                    <RANKING order="3" place="3" resultid="5114" />
                    <RANKING order="4" place="4" resultid="5508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1141" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5057" />
                    <RANKING order="2" place="2" resultid="5505" />
                    <RANKING order="3" place="3" resultid="5516" />
                    <RANKING order="4" place="4" resultid="5074" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1142" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5029" />
                    <RANKING order="2" place="2" resultid="5340" />
                    <RANKING order="3" place="3" resultid="5500" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4882" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4883" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4884" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4885" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1143" gender="F" number="19" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1144" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1145" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1146" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1147" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1148" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1149" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5050" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4886" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1151" gender="M" number="20" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1152" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5109" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1153" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1154" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5352" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1155" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1156" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5071" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1157" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1158" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4887" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1161" gender="M" number="22" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1162" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5470" />
                    <RANKING order="2" place="2" resultid="5289" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4888" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1163" gender="F" number="23" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1164" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5403" />
                    <RANKING order="2" place="2" resultid="5259" />
                    <RANKING order="3" place="3" resultid="5372" />
                    <RANKING order="4" place="4" resultid="5228" />
                    <RANKING order="5" place="5" resultid="5442" />
                    <RANKING order="6" place="6" resultid="5459" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1165" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5022" />
                    <RANKING order="2" place="2" resultid="5169" />
                    <RANKING order="3" place="3" resultid="5360" />
                    <RANKING order="4" place="4" resultid="5462" />
                    <RANKING order="5" place="5" resultid="5481" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4889" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4890" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1166" gender="M" number="24" order="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1167" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5301" />
                    <RANKING order="2" place="2" resultid="5256" />
                    <RANKING order="3" place="3" resultid="5024" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1168" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5223" />
                    <RANKING order="2" place="2" resultid="5305" />
                    <RANKING order="3" place="3" resultid="5280" />
                    <RANKING order="4" place="4" resultid="5318" />
                    <RANKING order="5" place="-1" resultid="5452" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4891" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4892" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1169" gender="F" number="25" order="23" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1170" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5395" />
                    <RANKING order="2" place="2" resultid="5207" />
                    <RANKING order="3" place="3" resultid="5368" />
                    <RANKING order="4" place="4" resultid="5411" />
                    <RANKING order="5" place="5" resultid="5422" />
                    <RANKING order="6" place="6" resultid="5268" />
                    <RANKING order="7" place="-1" resultid="5456" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1171" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5324" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4893" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4894" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1172" gender="M" number="26" order="24" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1173" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5153" />
                    <RANKING order="2" place="2" resultid="5314" />
                    <RANKING order="3" place="3" resultid="5449" />
                    <RANKING order="4" place="4" resultid="5138" />
                    <RANKING order="5" place="5" resultid="5379" />
                    <RANKING order="6" place="6" resultid="5297" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1174" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5202" />
                    <RANKING order="2" place="2" resultid="5127" />
                    <RANKING order="3" place="3" resultid="5474" />
                    <RANKING order="4" place="-1" resultid="5009" />
                    <RANKING order="5" place="-1" resultid="5484" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4895" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4896" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1175" gender="F" number="27" order="25" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1176" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1177" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1178" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5063" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1179" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1180" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5495" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1181" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1182" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5053" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4897" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1183" gender="M" number="28" order="26" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1184" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5383" />
                    <RANKING order="2" place="2" resultid="5119" />
                    <RANKING order="3" place="-1" resultid="5328" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1185" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5041" />
                    <RANKING order="2" place="2" resultid="5514" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5098" />
                    <RANKING order="2" place="2" resultid="5348" />
                    <RANKING order="3" place="3" resultid="5286" />
                    <RANKING order="4" place="4" resultid="5497" />
                    <RANKING order="5" place="5" resultid="5292" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1187" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4979" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1188" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1189" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5075" />
                    <RANKING order="2" place="2" resultid="5356" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1190" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5534" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4898" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4899" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4900" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1191" gender="F" number="29" order="27" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1192" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5344" />
                    <RANKING order="2" place="2" resultid="5237" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1193" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5083" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1194" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5093" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1195" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4991" />
                    <RANKING order="2" place="2" resultid="5332" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1196" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1197" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1198" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4901" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1199" gender="M" number="30" order="28" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1200" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1201" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5077" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1202" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1203" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1204" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1205" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1206" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5489" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4902" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2023-03-18" daytime="15:55" number="2" warmupfrom="14:45" warmupuntil="15:45">
          <EVENTS>
            <EVENT eventid="1207" gender="F" number="31" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1208" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5404" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1209" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5170" />
                    <RANKING order="2" place="2" resultid="5143" />
                    <RANKING order="3" place="3" resultid="5435" />
                    <RANKING order="4" place="4" resultid="5427" />
                    <RANKING order="5" place="5" resultid="5361" />
                    <RANKING order="6" place="6" resultid="5337" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4903" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4904" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1210" gender="M" number="32" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1211" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5302" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1212" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5181" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4905" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1213" gender="F" number="33" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1214" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4986" />
                    <RANKING order="2" place="2" resultid="5004" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1215" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1216" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5017" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1217" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4992" />
                    <RANKING order="2" place="2" resultid="5333" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1218" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1219" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1220" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4906" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1221" gender="M" number="34" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1222" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1223" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5078" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1224" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5032" />
                    <RANKING order="2" place="2" resultid="4998" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1225" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1226" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1227" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1228" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5341" />
                    <RANKING order="2" place="-1" resultid="5490" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4907" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1229" gender="F" number="35" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1230" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5412" />
                    <RANKING order="2" place="2" resultid="5431" />
                    <RANKING order="3" place="3" resultid="5365" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1231" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5148" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4908" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1232" gender="M" number="36" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1233" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5400" />
                    <RANKING order="2" place="2" resultid="5450" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1234" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5392" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4909" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1235" gender="F" number="37" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1236" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5345" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1237" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1238" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1239" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1240" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1241" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1242" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4910" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1243" gender="M" number="38" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1244" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5384" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1245" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5042" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1246" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5099" />
                    <RANKING order="2" place="2" resultid="5047" />
                    <RANKING order="3" place="3" resultid="5349" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1247" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4980" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1248" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1249" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5357" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1250" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5030" />
                    <RANKING order="2" place="-1" resultid="5535" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4911" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4912" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1253" gender="M" number="40" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1254" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5290" />
                    <RANKING order="2" place="2" resultid="5471" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4913" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1255" gender="F" number="41" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1256" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5229" />
                    <RANKING order="2" place="2" resultid="5373" />
                    <RANKING order="3" place="3" resultid="5443" />
                    <RANKING order="4" place="4" resultid="5260" />
                    <RANKING order="5" place="5" resultid="5531" />
                    <RANKING order="6" place="6" resultid="5466" />
                    <RANKING order="7" place="7" resultid="5460" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1257" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5023" />
                    <RANKING order="2" place="2" resultid="5338" />
                    <RANKING order="3" place="3" resultid="5428" />
                    <RANKING order="4" place="4" resultid="5171" />
                    <RANKING order="5" place="5" resultid="5144" />
                    <RANKING order="6" place="6" resultid="5463" />
                    <RANKING order="7" place="7" resultid="5376" />
                    <RANKING order="8" place="8" resultid="5482" />
                    <RANKING order="9" place="9" resultid="5213" />
                    <RANKING order="10" place="10" resultid="5362" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4914" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4915" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4916" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1258" gender="M" number="42" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1259" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5257" />
                    <RANKING order="2" place="2" resultid="5303" />
                    <RANKING order="3" place="3" resultid="5264" />
                    <RANKING order="4" place="4" resultid="5025" />
                    <RANKING order="5" place="5" resultid="5529" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1260" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5224" />
                    <RANKING order="2" place="2" resultid="5182" />
                    <RANKING order="3" place="3" resultid="5319" />
                    <RANKING order="4" place="4" resultid="5453" />
                    <RANKING order="5" place="5" resultid="5311" />
                    <RANKING order="6" place="6" resultid="5281" />
                    <RANKING order="7" place="7" resultid="5306" />
                    <RANKING order="8" place="8" resultid="5447" />
                    <RANKING order="9" place="9" resultid="5468" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4917" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4918" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4919" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1261" gender="F" number="43" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1262" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5423" />
                    <RANKING order="2" place="2" resultid="5208" />
                    <RANKING order="3" place="3" resultid="5218" />
                    <RANKING order="4" place="4" resultid="5369" />
                    <RANKING order="5" place="5" resultid="5408" />
                    <RANKING order="6" place="6" resultid="5165" />
                    <RANKING order="7" place="7" resultid="5366" />
                    <RANKING order="8" place="8" resultid="5527" />
                    <RANKING order="9" place="9" resultid="5523" />
                    <RANKING order="10" place="10" resultid="5253" />
                    <RANKING order="11" place="11" resultid="5457" />
                    <RANKING order="12" place="12" resultid="5269" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1263" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5133" />
                    <RANKING order="2" place="2" resultid="5149" />
                    <RANKING order="3" place="3" resultid="5277" />
                    <RANKING order="4" place="4" resultid="5325" />
                    <RANKING order="5" place="5" resultid="5284" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4920" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4921" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4922" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1264" gender="M" number="44" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1265" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5192" />
                    <RANKING order="2" place="2" resultid="5175" />
                    <RANKING order="3" place="3" resultid="5154" />
                    <RANKING order="4" place="4" resultid="5388" />
                    <RANKING order="5" place="5" resultid="5315" />
                    <RANKING order="6" place="6" resultid="5186" />
                    <RANKING order="7" place="7" resultid="5539" />
                    <RANKING order="8" place="8" resultid="5198" />
                    <RANKING order="9" place="9" resultid="5401" />
                    <RANKING order="10" place="10" resultid="5139" />
                    <RANKING order="11" place="11" resultid="5380" />
                    <RANKING order="12" place="12" resultid="5525" />
                    <RANKING order="13" place="13" resultid="5298" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1266" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5416" />
                    <RANKING order="2" place="2" resultid="5203" />
                    <RANKING order="3" place="3" resultid="5393" />
                    <RANKING order="4" place="4" resultid="5128" />
                    <RANKING order="5" place="5" resultid="5010" />
                    <RANKING order="6" place="6" resultid="5439" />
                    <RANKING order="7" place="7" resultid="5475" />
                    <RANKING order="8" place="8" resultid="5273" />
                    <RANKING order="9" place="9" resultid="5533" />
                    <RANKING order="10" place="10" resultid="5485" />
                    <RANKING order="11" place="11" resultid="5488" />
                    <RANKING order="12" place="-1" resultid="5124" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4923" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4924" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4925" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4926" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1267" gender="F" number="45" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1268" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5243" />
                    <RANKING order="2" place="2" resultid="4987" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1269" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5088" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1270" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5094" />
                    <RANKING order="2" place="2" resultid="5064" />
                    <RANKING order="3" place="3" resultid="5018" />
                    <RANKING order="4" place="4" resultid="5248" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1271" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1272" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5496" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1273" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5059" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1274" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4927" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4928" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1275" gender="M" number="46" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1276" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5120" />
                    <RANKING order="2" place="2" resultid="5329" />
                    <RANKING order="3" place="3" resultid="5385" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1277" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5104" />
                    <RANKING order="2" place="2" resultid="5515" />
                    <RANKING order="3" place="3" resultid="5419" />
                    <RANKING order="4" place="4" resultid="5159" />
                    <RANKING order="5" place="-1" resultid="5503" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1278" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5033" />
                    <RANKING order="2" place="2" resultid="5037" />
                    <RANKING order="3" place="3" resultid="5353" />
                    <RANKING order="4" place="4" resultid="5498" />
                    <RANKING order="5" place="5" resultid="5287" />
                    <RANKING order="6" place="6" resultid="5293" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1279" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5512" />
                    <RANKING order="2" place="2" resultid="5520" />
                    <RANKING order="3" place="3" resultid="5234" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1280" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5027" />
                    <RANKING order="2" place="2" resultid="5115" />
                    <RANKING order="3" place="3" resultid="5509" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1281" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5506" />
                    <RANKING order="2" place="2" resultid="5517" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1282" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5492" />
                    <RANKING order="2" place="2" resultid="5321" />
                    <RANKING order="3" place="3" resultid="5501" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4929" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4930" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4931" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4932" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1283" gender="F" number="47" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1284" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5238" />
                    <RANKING order="2" place="-1" resultid="5005" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1285" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5084" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1286" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1287" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5334" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1288" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1289" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1290" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4933" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1291" gender="M" number="48" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1292" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5110" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1293" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5420" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1294" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4999" />
                    <RANKING order="2" place="2" resultid="5068" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1295" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1296" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1297" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1298" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="5342" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4934" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1301" gender="M" number="50" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1302" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5472" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4935" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1303" gender="F" number="51" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1304" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5405" />
                    <RANKING order="2" place="2" resultid="5230" />
                    <RANKING order="3" place="3" resultid="5261" />
                    <RANKING order="4" place="4" resultid="5444" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1305" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5436" />
                    <RANKING order="2" place="2" resultid="5464" />
                    <RANKING order="3" place="3" resultid="5377" />
                    <RANKING order="4" place="4" resultid="5214" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4936" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4937" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1306" gender="M" number="52" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1307" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5258" />
                    <RANKING order="2" place="2" resultid="5265" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1308" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5225" />
                    <RANKING order="2" place="2" resultid="5312" />
                    <RANKING order="3" place="3" resultid="5320" />
                    <RANKING order="4" place="4" resultid="5307" />
                    <RANKING order="5" place="5" resultid="5282" />
                    <RANKING order="6" place="-1" resultid="5454" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4938" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4939" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1309" gender="F" number="53" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1310" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5396" />
                    <RANKING order="2" place="2" resultid="5409" />
                    <RANKING order="3" place="3" resultid="5432" />
                    <RANKING order="4" place="4" resultid="5219" />
                    <RANKING order="5" place="5" resultid="5254" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1311" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5134" />
                    <RANKING order="2" place="2" resultid="5278" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4940" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4941" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1312" gender="M" number="54" order="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1313" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5193" />
                    <RANKING order="2" place="2" resultid="5155" />
                    <RANKING order="3" place="3" resultid="5176" />
                    <RANKING order="4" place="4" resultid="5389" />
                    <RANKING order="5" place="5" resultid="5187" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1314" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5440" />
                    <RANKING order="2" place="2" resultid="5478" />
                    <RANKING order="3" place="-1" resultid="5125" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4942" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4943" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1315" gender="F" number="55" order="23" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1316" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5244" />
                    <RANKING order="2" place="2" resultid="5346" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1317" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5089" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1318" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5095" />
                    <RANKING order="2" place="2" resultid="5065" />
                    <RANKING order="3" place="3" resultid="5249" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1319" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1320" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1321" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1322" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4944" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1323" gender="M" number="56" order="24" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1324" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5330" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1325" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5105" />
                    <RANKING order="2" place="2" resultid="5043" />
                    <RANKING order="3" place="3" resultid="5160" />
                    <RANKING order="4" place="-1" resultid="5504" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1326" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5354" />
                    <RANKING order="2" place="2" resultid="5038" />
                    <RANKING order="3" place="3" resultid="5294" />
                    <RANKING order="4" place="-1" resultid="5499" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1327" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4981" />
                    <RANKING order="2" place="2" resultid="5521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1328" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5510" />
                    <RANKING order="2" place="2" resultid="5116" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1329" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5507" />
                    <RANKING order="2" place="2" resultid="5518" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1330" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5493" />
                    <RANKING order="2" place="2" resultid="5322" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4945" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4946" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4947" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1331" gender="F" number="57" order="25" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1332" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1333" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1334" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1335" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1336" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1337" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1338" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5054" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4948" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1339" gender="M" number="58" order="26" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1340" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="5111" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1341" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5079" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1342" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5048" />
                    <RANKING order="2" place="2" resultid="5350" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1343" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1344" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5072" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1345" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5358" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1346" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4949" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1347" gender="F" number="59" order="27" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1348" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5397" />
                    <RANKING order="2" place="2" resultid="5413" />
                    <RANKING order="3" place="3" resultid="5209" />
                    <RANKING order="4" place="4" resultid="5370" />
                    <RANKING order="5" place="5" resultid="5424" />
                    <RANKING order="6" place="6" resultid="5270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1349" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5326" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4950" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4951" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1350" gender="M" number="60" order="28" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1351" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5316" />
                    <RANKING order="2" place="2" resultid="5451" />
                    <RANKING order="3" place="3" resultid="5140" />
                    <RANKING order="4" place="4" resultid="5381" />
                    <RANKING order="5" place="5" resultid="5299" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1352" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5204" />
                    <RANKING order="2" place="2" resultid="5129" />
                    <RANKING order="3" place="3" resultid="5011" />
                    <RANKING order="4" place="-1" resultid="5479" />
                    <RANKING order="5" place="-1" resultid="5486" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4952" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4953" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2023-03-19" daytime="09:10" number="3" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="1353" gender="F" number="61" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1354" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5245" />
                    <RANKING order="2" place="2" resultid="4988" />
                    <RANKING order="3" place="3" resultid="5239" />
                    <RANKING order="4" place="4" resultid="5006" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1355" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5090" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1356" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5066" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1357" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4994" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1358" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1359" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1360" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4954" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4955" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1361" gender="M" number="62" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1362" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5112" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1363" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5080" />
                    <RANKING order="2" place="2" resultid="5106" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1364" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5034" />
                    <RANKING order="2" place="2" resultid="5039" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1365" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5235" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1366" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5028" />
                    <RANKING order="2" place="2" resultid="5117" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1367" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5519" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1368" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4956" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4957" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1369" gender="F" number="63" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1370" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1371" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1372" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5019" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1373" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1374" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1375" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1376" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5055" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4958" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1377" gender="M" number="64" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1378" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1379" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5044" />
                    <RANKING order="2" place="2" resultid="5161" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1380" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5100" />
                    <RANKING order="2" place="2" resultid="5049" />
                    <RANKING order="3" place="3" resultid="5295" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1381" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4982" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1382" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1383" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1384" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5536" />
                    <RANKING order="2" place="2" resultid="5502" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4959" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4960" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1389" gender="F" number="67" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1390" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="5166" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1391" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5150" />
                    <RANKING order="2" place="2" resultid="5013" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4961" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1392" gender="M" number="68" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1393" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5194" />
                    <RANKING order="2" place="2" resultid="5177" />
                    <RANKING order="3" place="3" resultid="5199" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1394" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="5274" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4962" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1395" gender="F" number="69" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1396" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5240" />
                    <RANKING order="2" place="2" resultid="4989" />
                    <RANKING order="3" place="3" resultid="5007" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1397" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5085" />
                    <RANKING order="2" place="2" resultid="5091" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1398" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1399" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1400" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1401" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1402" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4963" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1403" gender="M" number="70" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1404" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5121" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1405" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1406" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5101" />
                    <RANKING order="2" place="2" resultid="5000" />
                    <RANKING order="3" place="3" resultid="5040" />
                    <RANKING order="4" place="4" resultid="5069" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1407" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1408" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1409" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1410" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4964" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1411" gender="F" number="71" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1412" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5231" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1413" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5145" />
                    <RANKING order="2" place="2" resultid="5172" />
                    <RANKING order="3" place="3" resultid="5215" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4965" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1414" gender="M" number="72" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1415" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5266" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1416" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5226" />
                    <RANKING order="2" place="2" resultid="5183" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4966" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1417" gender="F" number="73" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1418" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5210" />
                    <RANKING order="2" place="2" resultid="5220" />
                    <RANKING order="3" place="3" resultid="5167" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1419" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5135" />
                    <RANKING order="2" place="2" resultid="5151" />
                    <RANKING order="3" place="3" resultid="5014" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4967" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1420" gender="M" number="74" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1421" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5195" />
                    <RANKING order="2" place="2" resultid="5178" />
                    <RANKING order="3" place="3" resultid="5156" />
                    <RANKING order="4" place="4" resultid="5200" />
                    <RANKING order="5" place="5" resultid="5188" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1422" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5130" />
                    <RANKING order="2" place="2" resultid="5205" />
                    <RANKING order="3" place="3" resultid="5012" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4968" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4969" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1423" gender="F" number="75" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1424" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1425" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5086" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1426" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5020" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1427" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1428" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1429" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1430" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4970" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1431" gender="M" number="76" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1432" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1433" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5045" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1434" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1435" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1436" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1437" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1438" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4971" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1439" gender="F" number="77" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1440" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="5221" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1441" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5136" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4972" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1442" gender="M" number="78" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1443" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5189" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1444" agemax="12" agemin="12" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4973" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1445" gender="F" number="79" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1446" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5246" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1447" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1448" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5096" />
                    <RANKING order="2" place="2" resultid="5250" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1449" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4995" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1450" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1451" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5051" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1452" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4974" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1453" gender="M" number="80" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1454" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5113" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1455" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5107" />
                    <RANKING order="2" place="-1" resultid="5162" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1456" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5035" />
                    <RANKING order="2" place="2" resultid="5001" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1457" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4983" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1458" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5073" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1459" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1460" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4975" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4976" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1469" gender="M" number="82" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1470" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1471" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5081" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1472" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1473" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1474" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1475" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1476" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4977" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="16053" nation="BRA" clubid="4576" swrid="93777" name="Fábrica de Nadadores" shortname="Fábrica">
          <ATHLETES>
            <ATHLETE firstname="Kenzo" lastname="Toshiro Miura" birthdate="2011-04-05" gender="M" nation="BRA" license="391850" swrid="5603921" athleteid="4761" externalid="391850">
              <RESULTS>
                <RESULT eventid="1096" points="101" reactiontime="0" swimtime="00:00:47.63" resultid="5476" heatid="4863" lane="3" />
                <RESULT eventid="1124" points="102" reactiontime="0" swimtime="00:01:35.87" resultid="5477" heatid="4876" lane="3" />
                <RESULT eventid="1312" points="66" reactiontime="0" swimtime="00:00:53.81" resultid="5478" heatid="4942" lane="3" />
                <RESULT eventid="1350" reactiontime="0" status="DSQ" swimtime="00:00:00.00" resultid="5479" heatid="4952" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabel" lastname="Rezende" birthdate="2013-12-13" gender="F" nation="BRA" license="370657" swrid="5603900" athleteid="4587" externalid="370657">
              <RESULTS>
                <RESULT eventid="1087" points="116" reactiontime="0" swimtime="00:00:51.71" resultid="5335" heatid="4859" lane="6" entrytime="00:00:59.03" />
                <RESULT eventid="1115" points="110" reactiontime="0" swimtime="00:01:44.65" resultid="5336" heatid="4871" lane="6" entrytime="00:01:54.14" />
                <RESULT eventid="1207" points="81" reactiontime="0" swimtime="00:02:10.17" resultid="5337" heatid="4904" lane="5" entrytime="00:02:45.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1255" points="139" reactiontime="0" swimtime="00:00:44.20" resultid="5338" heatid="4916" lane="6" entrytime="00:00:50.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alex" lastname="Junior" birthdate="2013-03-11" gender="M" nation="BRA" license="385710" swrid="5603860" athleteid="4720" externalid="385710">
              <RESULTS>
                <RESULT eventid="1090" points="37" reactiontime="0" swimtime="00:01:06.20" resultid="5445" heatid="4860" lane="5" entrytime="00:01:31.35" />
                <RESULT eventid="1118" points="20" reactiontime="0" swimtime="00:02:43.17" resultid="5446" heatid="4872" lane="4" />
                <RESULT eventid="1258" points="38" reactiontime="0" swimtime="00:00:59.91" resultid="5447" heatid="4919" lane="3" entrytime="00:01:19.36" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Gabriel Ribeiro" birthdate="2011-06-23" gender="M" nation="BRA" license="392052" swrid="5603839" athleteid="4770" externalid="392052">
              <RESULTS>
                <RESULT eventid="1124" points="46" reactiontime="0" swimtime="00:02:04.90" resultid="5483" heatid="4877" lane="3" />
                <RESULT eventid="1172" reactiontime="0" status="DNS" swimtime="00:00:00.00" resultid="5484" />
                <RESULT eventid="1264" points="59" reactiontime="0" swimtime="00:00:51.63" resultid="5485" heatid="4924" lane="2" />
                <RESULT eventid="1350" reactiontime="0" status="DSQ" swimtime="00:00:00.00" resultid="5486" heatid="4953" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Bertão" birthdate="2012-05-23" gender="M" nation="BRA" license="378344" swrid="5306272" athleteid="4636" externalid="378344">
              <RESULTS>
                <RESULT eventid="1124" points="48" reactiontime="0" swimtime="00:02:03.35" resultid="5378" heatid="4877" lane="5" entrytime="00:02:11.31" />
                <RESULT eventid="1172" points="57" reactiontime="0" swimtime="00:01:04.48" resultid="5379" heatid="4895" lane="4" entrytime="00:01:04.79" />
                <RESULT eventid="1264" points="48" reactiontime="0" swimtime="00:00:55.38" resultid="5380" heatid="4924" lane="5" entrytime="00:00:59.16" />
                <RESULT eventid="1350" points="52" reactiontime="0" swimtime="00:02:27.47" resultid="5381" heatid="4952" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Perola" lastname="Maria Hamerschimidt" birthdate="2014-08-20" gender="F" nation="BRA" license="391846" swrid="5603868" athleteid="4746" externalid="391846">
              <RESULTS>
                <RESULT eventid="1087" points="28" reactiontime="0" swimtime="00:01:23.21" resultid="5465" heatid="4858" lane="6" />
                <RESULT eventid="1255" points="35" reactiontime="0" swimtime="00:01:09.97" resultid="5466" heatid="4914" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Tiemi Yamaguchi" birthdate="2013-02-28" gender="F" nation="BRA" license="385707" swrid="5603920" athleteid="4705" externalid="385707">
              <RESULTS>
                <RESULT eventid="1087" points="113" reactiontime="0" swimtime="00:00:52.14" resultid="5433" heatid="4859" lane="2" entrytime="00:01:02.09" />
                <RESULT eventid="1115" points="106" reactiontime="0" swimtime="00:01:45.89" resultid="5434" heatid="4871" lane="3" entrytime="00:01:50.85" />
                <RESULT eventid="1207" points="118" reactiontime="0" swimtime="00:01:55.21" resultid="5435" heatid="4903" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1303" points="102" reactiontime="0" swimtime="00:00:52.08" resultid="5436" heatid="4937" lane="6" entrytime="00:01:12.04" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Bagatim" birthdate="2014-05-27" gender="F" nation="BRA" license="378353" swrid="5236649" athleteid="4666" externalid="378353">
              <RESULTS>
                <RESULT eventid="1115" points="152" reactiontime="0" swimtime="00:01:34.00" resultid="5402" heatid="4869" lane="3" />
                <RESULT eventid="1163" points="146" reactiontime="0" swimtime="00:00:54.13" resultid="5403" heatid="4890" lane="4" entrytime="00:00:52.39" />
                <RESULT eventid="1207" points="140" reactiontime="0" swimtime="00:01:48.60" resultid="5404" heatid="4904" lane="6" />
                <RESULT eventid="1303" points="119" reactiontime="0" swimtime="00:00:49.45" resultid="5405" heatid="4937" lane="4" entrytime="00:00:46.26" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tiago" lastname="Mesti Bonetti" birthdate="2011-11-21" gender="M" nation="BRA" license="391849" swrid="5603874" athleteid="4757" externalid="391849">
              <RESULTS>
                <RESULT eventid="1124" points="63" reactiontime="0" swimtime="00:01:52.15" resultid="5473" heatid="4877" lane="6" />
                <RESULT eventid="1172" points="67" reactiontime="0" swimtime="00:01:01.18" resultid="5474" heatid="4895" lane="5" />
                <RESULT eventid="1264" points="102" reactiontime="0" swimtime="00:00:43.07" resultid="5475" heatid="4923" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monique" lastname="Istake" birthdate="2012-04-03" gender="F" nation="BRA" license="372023" swrid="5603857" athleteid="4676" externalid="372023">
              <RESULTS>
                <RESULT eventid="1061" points="196" reactiontime="0" swimtime="00:03:29.56" resultid="5410" heatid="4851" lane="6" entrytime="00:04:04.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.24" />
                    <SPLIT distance="100" swimtime="00:01:39.20" />
                    <SPLIT distance="150" swimtime="00:02:44.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1169" points="191" reactiontime="0" swimtime="00:00:49.51" resultid="5411" heatid="4893" lane="4" entrytime="00:01:12.28" />
                <RESULT eventid="1229" points="225" reactiontime="0" swimtime="00:06:24.32" resultid="5412" heatid="4908" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.62" />
                    <SPLIT distance="100" swimtime="00:01:31.62" />
                    <SPLIT distance="150" swimtime="00:02:20.81" />
                    <SPLIT distance="200" swimtime="00:03:09.40" />
                    <SPLIT distance="250" swimtime="00:03:59.48" />
                    <SPLIT distance="300" swimtime="00:04:48.85" />
                    <SPLIT distance="350" swimtime="00:05:38.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1347" points="183" reactiontime="0" swimtime="00:01:49.77" resultid="5413" heatid="4950" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Mendes Costa" birthdate="2014-04-03" gender="F" nation="BRA" license="378341" swrid="5603873" athleteid="4627" externalid="378341">
              <RESULTS>
                <RESULT eventid="1115" points="77" reactiontime="0" swimtime="00:01:58.08" resultid="5371" heatid="4870" lane="3" />
                <RESULT eventid="1163" points="77" reactiontime="0" swimtime="00:01:06.90" resultid="5372" heatid="4889" lane="2" />
                <RESULT eventid="1255" points="84" reactiontime="0" swimtime="00:00:52.19" resultid="5373" heatid="4914" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Guinoza" birthdate="2013-01-06" gender="F" nation="BRA" license="392012" swrid="5510698" athleteid="4766" externalid="392012">
              <RESULTS>
                <RESULT eventid="1115" points="99" reactiontime="0" swimtime="00:01:48.29" resultid="5480" heatid="4869" lane="5" />
                <RESULT eventid="1163" points="65" reactiontime="0" swimtime="00:01:10.95" resultid="5481" heatid="4890" lane="2" />
                <RESULT eventid="1255" points="101" reactiontime="0" swimtime="00:00:49.13" resultid="5482" heatid="4914" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Guilherme Ortega" birthdate="1999-08-05" gender="M" nation="BRA" license="383118" swrid="5603852" athleteid="4582" externalid="383118">
              <RESULTS>
                <RESULT eventid="1107" points="304" reactiontime="0" swimtime="00:00:33.03" resultid="5339" heatid="4868" lane="5" entrytime="00:00:32.49" />
                <RESULT eventid="1135" points="298" reactiontime="0" swimtime="00:01:07.13" resultid="5340" heatid="4882" lane="3" />
                <RESULT eventid="1221" points="221" reactiontime="0" swimtime="00:05:50.94" resultid="5341" heatid="4907" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                    <SPLIT distance="100" swimtime="00:01:14.14" />
                    <SPLIT distance="150" swimtime="00:01:58.22" />
                    <SPLIT distance="200" swimtime="00:02:43.28" />
                    <SPLIT distance="250" swimtime="00:03:29.81" />
                    <SPLIT distance="300" swimtime="00:04:17.12" />
                    <SPLIT distance="350" swimtime="00:05:05.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1291" reactiontime="0" status="DSQ" swimtime="00:00:00.00" resultid="5342" heatid="4934" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.42" />
                    <SPLIT distance="100" swimtime="00:01:19.52" />
                    <SPLIT distance="150" swimtime="00:02:03.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andressa" lastname="Zamarian Gouvea" birthdate="2007-09-18" gender="F" nation="BRA" license="318503" swrid="5603929" athleteid="4577" externalid="318503">
              <RESULTS>
                <RESULT eventid="1099" points="367" reactiontime="0" swimtime="00:00:35.29" resultid="5331" heatid="4866" lane="4" entrytime="00:00:36.53" />
                <RESULT eventid="1191" points="378" reactiontime="0" swimtime="00:11:02.38" resultid="5332" heatid="4901" lane="3" entrytime="00:10:59.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:11:04.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="382" reactiontime="0" swimtime="00:05:22.26" resultid="5333" heatid="4906" lane="5" entrytime="00:05:16.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                    <SPLIT distance="100" swimtime="00:01:14.44" />
                    <SPLIT distance="150" swimtime="00:01:56.29" />
                    <SPLIT distance="200" swimtime="00:02:37.79" />
                    <SPLIT distance="250" swimtime="00:03:20.17" />
                    <SPLIT distance="300" swimtime="00:04:03.14" />
                    <SPLIT distance="350" swimtime="00:04:44.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1283" points="350" reactiontime="0" swimtime="00:02:48.75" resultid="5334" heatid="4933" lane="4" entrytime="00:02:43.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.45" />
                    <SPLIT distance="100" swimtime="00:01:21.50" />
                    <SPLIT distance="150" swimtime="00:02:08.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruna" lastname="Scalise Drapzichinski" birthdate="2012-03-07" gender="F" nation="BRA" license="378349" swrid="5603909" athleteid="4656" externalid="378349">
              <RESULTS>
                <RESULT eventid="1061" points="208" reactiontime="0" swimtime="00:03:25.60" resultid="5394" heatid="4851" lane="5" entrytime="00:03:44.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.55" />
                    <SPLIT distance="100" swimtime="00:01:40.14" />
                    <SPLIT distance="150" swimtime="00:02:39.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1169" points="260" reactiontime="0" swimtime="00:00:44.70" resultid="5395" heatid="4894" lane="4" entrytime="00:00:50.06" />
                <RESULT eventid="1309" points="170" reactiontime="0" swimtime="00:00:43.96" resultid="5396" heatid="4940" lane="4" />
                <RESULT eventid="1347" points="222" reactiontime="0" swimtime="00:01:42.89" resultid="5397" heatid="4951" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eloah" lastname="Frasson" birthdate="2012-06-14" gender="F" nation="BRA" license="378338" swrid="5577016" athleteid="4622" externalid="378338">
              <RESULTS>
                <RESULT eventid="1121" points="132" reactiontime="0" swimtime="00:01:38.56" resultid="5367" heatid="4875" lane="6" entrytime="00:01:48.70" />
                <RESULT eventid="1169" points="197" reactiontime="0" swimtime="00:00:49.03" resultid="5368" heatid="4894" lane="6" entrytime="00:00:54.24" />
                <RESULT eventid="1261" points="163" reactiontime="0" swimtime="00:00:41.92" resultid="5369" heatid="4921" lane="4" entrytime="00:00:50.17" />
                <RESULT eventid="1347" points="172" reactiontime="0" swimtime="00:01:52.09" resultid="5370" heatid="4951" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vittorio" lastname="Furquim Marson" birthdate="2013-05-10" gender="M" nation="BRA" license="391842" swrid="5601999" athleteid="4729" externalid="391842">
              <RESULTS>
                <RESULT eventid="1166" reactiontime="0" status="DNS" swimtime="00:00:00.00" resultid="5452" />
                <RESULT eventid="1258" points="82" reactiontime="0" swimtime="00:00:46.38" resultid="5453" heatid="4918" lane="5" />
                <RESULT eventid="1306" reactiontime="0" status="DNS" swimtime="00:00:00.00" resultid="5454" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Braga" birthdate="2010-05-07" gender="M" nation="BRA" license="378345" swrid="5343953" athleteid="4641" externalid="378345">
              <RESULTS>
                <RESULT eventid="1075" points="193" reactiontime="0" swimtime="00:03:09.55" resultid="5382" heatid="4854" lane="5" />
                <RESULT eventid="1183" points="221" reactiontime="0" swimtime="00:00:41.24" resultid="5383" heatid="4899" lane="4" entrytime="00:00:43.81" />
                <RESULT eventid="1243" points="231" reactiontime="0" swimtime="00:03:15.61" resultid="5384" heatid="4911" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.25" />
                    <SPLIT distance="100" swimtime="00:01:33.13" />
                    <SPLIT distance="150" swimtime="00:02:25.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1275" points="160" reactiontime="0" swimtime="00:00:37.08" resultid="5385" heatid="4929" lane="4" entrytime="00:00:38.89" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Gevaerd Verssutti Garcia" birthdate="2013-10-15" gender="F" nation="BRA" license="378404" swrid="5588723" athleteid="4695" externalid="378404">
              <RESULTS>
                <RESULT eventid="1087" points="143" reactiontime="0" swimtime="00:00:48.23" resultid="5425" heatid="4859" lane="4" entrytime="00:00:50.68" />
                <RESULT eventid="1115" points="131" reactiontime="0" swimtime="00:01:38.74" resultid="5426" heatid="4871" lane="4" entrytime="00:01:41.45" />
                <RESULT eventid="1207" points="109" reactiontime="0" swimtime="00:01:57.94" resultid="5427" heatid="4903" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1255" points="137" reactiontime="0" swimtime="00:00:44.44" resultid="5428" heatid="4916" lane="5" entrytime="00:00:40.92" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Sachetti Fabian" birthdate="2012-08-09" gender="F" nation="BRA" license="391843" swrid="5603903" athleteid="4733" externalid="391843">
              <RESULTS>
                <RESULT eventid="1093" points="68" reactiontime="0" swimtime="00:01:01.74" resultid="5455" heatid="4861" lane="5" />
                <RESULT eventid="1169" reactiontime="0" status="DNS" swimtime="00:00:00.00" resultid="5456" />
                <RESULT eventid="1261" points="51" reactiontime="0" swimtime="00:01:01.72" resultid="5457" heatid="4920" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Jupi Takaki" birthdate="2013-03-26" gender="F" nation="BRA" license="391845" swrid="5603861" athleteid="4741" externalid="391845">
              <RESULTS>
                <RESULT eventid="1115" points="98" reactiontime="0" swimtime="00:01:48.76" resultid="5461" heatid="4869" lane="4" />
                <RESULT eventid="1163" points="76" reactiontime="0" swimtime="00:01:07.32" resultid="5462" heatid="4889" lane="5" />
                <RESULT eventid="1255" points="129" reactiontime="0" swimtime="00:00:45.37" resultid="5463" heatid="4915" lane="2" />
                <RESULT eventid="1303" points="82" reactiontime="0" swimtime="00:00:56.10" resultid="5464" heatid="4936" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amanda" lastname="Guerra" birthdate="2013-11-22" gender="F" nation="BRA" license="378336" swrid="5603849" athleteid="4612" externalid="378336">
              <RESULTS>
                <RESULT eventid="1115" points="79" reactiontime="0" swimtime="00:01:57.09" resultid="5359" heatid="4870" lane="6" />
                <RESULT eventid="1163" points="83" reactiontime="0" swimtime="00:01:05.30" resultid="5360" heatid="4889" lane="6" />
                <RESULT eventid="1207" points="84" reactiontime="0" swimtime="00:02:08.53" resultid="5361" heatid="4903" lane="5" />
                <RESULT eventid="1255" points="71" reactiontime="0" swimtime="00:00:55.13" resultid="5362" heatid="4915" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Pazinato" birthdate="2011-01-05" gender="M" nation="BRA" license="368149" swrid="5603889" athleteid="4681" externalid="368149">
              <RESULTS>
                <RESULT eventid="1096" points="164" reactiontime="0" swimtime="00:00:40.54" resultid="5414" heatid="4865" lane="3" entrytime="00:00:46.59" />
                <RESULT eventid="1124" points="204" reactiontime="0" swimtime="00:01:16.05" resultid="5415" heatid="4879" lane="5" entrytime="00:01:18.99" />
                <RESULT eventid="1264" points="200" reactiontime="0" swimtime="00:00:34.47" resultid="5416" heatid="4926" lane="4" entrytime="00:00:34.98" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Silveira De Almeida" birthdate="2008-07-08" gender="M" nation="BRA" license="368152" swrid="5603912" athleteid="4602" externalid="368152">
              <RESULTS>
                <RESULT eventid="1107" points="255" reactiontime="0" swimtime="00:00:35.02" resultid="5351" heatid="4868" lane="2" entrytime="00:00:47.06" />
                <RESULT eventid="1151" points="402" reactiontime="0" swimtime="00:02:26.63" resultid="5352" heatid="4887" lane="5" entrytime="00:03:14.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                    <SPLIT distance="100" swimtime="00:01:12.52" />
                    <SPLIT distance="150" swimtime="00:01:50.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1275" points="284" reactiontime="0" swimtime="00:00:30.64" resultid="5353" heatid="4931" lane="7" entrytime="00:00:32.98" />
                <RESULT eventid="1323" points="300" reactiontime="0" swimtime="00:00:32.49" resultid="5354" heatid="4947" lane="5" entrytime="00:00:30.58" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Silverio Duarte" birthdate="2011-08-08" gender="M" nation="BRA" license="392138" swrid="5603913" athleteid="4775" externalid="392138">
              <RESULTS>
                <RESULT eventid="1096" reactiontime="0" status="DSQ" swimtime="00:00:00.00" resultid="5487" heatid="4864" lane="2" />
                <RESULT eventid="1264" points="36" reactiontime="0" swimtime="00:01:00.65" resultid="5488" heatid="4923" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Valentina Gozaga" birthdate="2014-06-28" gender="F" nation="BRA" license="385709" swrid="5603924" athleteid="4715" externalid="385709">
              <RESULTS>
                <RESULT eventid="1115" points="70" reactiontime="0" swimtime="00:02:01.59" resultid="5441" heatid="4870" lane="4" />
                <RESULT eventid="1163" points="49" reactiontime="0" swimtime="00:01:18.02" resultid="5442" heatid="4890" lane="3" entrytime="00:01:22.46" />
                <RESULT eventid="1255" points="68" reactiontime="0" swimtime="00:00:55.94" resultid="5443" heatid="4916" lane="7" entrytime="00:00:54.84" />
                <RESULT eventid="1303" points="35" reactiontime="0" swimtime="00:01:14.51" resultid="5444" heatid="4937" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Posser" birthdate="2013-02-07" gender="F" nation="BRA" license="378343" swrid="5603896" athleteid="4631" externalid="378343">
              <RESULTS>
                <RESULT eventid="1087" points="84" reactiontime="0" swimtime="00:00:57.53" resultid="5374" heatid="4858" lane="4" entrytime="00:01:13.21" />
                <RESULT eventid="1115" points="77" reactiontime="0" swimtime="00:01:58.03" resultid="5375" heatid="4871" lane="7" entrytime="00:02:14.23" />
                <RESULT eventid="1255" points="126" reactiontime="0" swimtime="00:00:45.69" resultid="5376" heatid="4915" lane="4" entrytime="00:01:00.08" />
                <RESULT eventid="1303" points="65" reactiontime="0" swimtime="00:01:00.39" resultid="5377" heatid="4937" lane="5" entrytime="00:01:07.79" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="Sabaini Preis" birthdate="2013-08-20" gender="M" nation="BRA" license="391847" swrid="5603902" athleteid="4749" externalid="391847">
              <RESULTS>
                <RESULT eventid="1090" points="31" reactiontime="0" swimtime="00:01:10.40" resultid="5467" heatid="4860" lane="2" />
                <RESULT eventid="1258" points="28" reactiontime="0" swimtime="00:01:05.81" resultid="5468" heatid="4918" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bárbara" lastname="Maria Barreto" birthdate="2012-10-25" gender="F" nation="BRA" license="370672" swrid="5603867" athleteid="4671" externalid="370672">
              <RESULTS>
                <RESULT eventid="1093" points="123" reactiontime="0" swimtime="00:00:50.71" resultid="5406" heatid="4862" lane="5" entrytime="00:00:51.15" />
                <RESULT eventid="1061" points="156" reactiontime="0" swimtime="00:03:46.23" resultid="5407" heatid="4850" lane="4" />
                <RESULT eventid="1261" points="160" reactiontime="0" swimtime="00:00:42.17" resultid="5408" heatid="4922" lane="6" entrytime="00:00:43.74" />
                <RESULT eventid="1309" points="120" reactiontime="0" swimtime="00:00:49.38" resultid="5409" heatid="4941" lane="5" entrytime="00:00:59.68" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Kenji Yamaguchi" birthdate="2011-08-25" gender="M" nation="BRA" license="385708" swrid="5603862" athleteid="4710" externalid="385708">
              <RESULTS>
                <RESULT eventid="1064" points="123" reactiontime="0" swimtime="00:03:40.27" resultid="5437" heatid="4852" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.03" />
                    <SPLIT distance="100" swimtime="00:01:44.29" />
                    <SPLIT distance="150" swimtime="00:02:49.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="145" reactiontime="0" swimtime="00:01:25.28" resultid="5438" heatid="4878" lane="2" entrytime="00:01:47.94" />
                <RESULT eventid="1264" points="125" reactiontime="0" swimtime="00:00:40.30" resultid="5439" heatid="4924" lane="3" entrytime="00:01:00.15" />
                <RESULT eventid="1312" points="101" reactiontime="0" swimtime="00:00:46.65" resultid="5440" heatid="4943" lane="3" entrytime="00:00:49.51" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Drapzichinski" birthdate="2015-08-21" gender="M" nation="BRA" license="391848" swrid="5603890" athleteid="4752" externalid="391848">
              <RESULTS>
                <RESULT eventid="1085" points="50" reactiontime="0" swimtime="00:00:28.04" resultid="5469" heatid="4857" lane="4" />
                <RESULT eventid="1161" points="35" reactiontime="0" swimtime="00:00:35.04" resultid="5470" heatid="4888" lane="4" />
                <RESULT eventid="1253" points="29" reactiontime="0" swimtime="00:00:29.28" resultid="5471" heatid="4913" lane="4" />
                <RESULT eventid="1301" points="23" reactiontime="0" swimtime="00:00:34.30" resultid="5472" heatid="4935" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Sachetti Fabian" birthdate="2014-08-02" gender="F" nation="BRA" license="391844" swrid="5603904" athleteid="4737" externalid="391844">
              <RESULTS>
                <RESULT eventid="1087" points="37" reactiontime="0" swimtime="00:01:15.58" resultid="5458" heatid="4858" lane="3" />
                <RESULT eventid="1163" points="47" reactiontime="0" swimtime="00:01:18.91" resultid="5459" heatid="4890" lane="6" />
                <RESULT eventid="1255" points="20" reactiontime="0" swimtime="00:01:24.03" resultid="5460" heatid="4914" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Berto" birthdate="2008-10-22" gender="M" nation="BRA" license="378342" swrid="5312223" athleteid="4597" externalid="378342">
              <RESULTS>
                <RESULT eventid="1107" points="151" reactiontime="0" swimtime="00:00:41.65" resultid="5347" heatid="4867" lane="4" />
                <RESULT eventid="1183" points="253" reactiontime="0" swimtime="00:00:39.43" resultid="5348" heatid="4900" lane="7" entrytime="00:00:41.97" />
                <RESULT eventid="1243" points="286" reactiontime="0" swimtime="00:03:02.34" resultid="5349" heatid="4911" lane="4" entrytime="00:03:04.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.30" />
                    <SPLIT distance="100" swimtime="00:01:26.56" />
                    <SPLIT distance="150" swimtime="00:02:14.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1339" points="210" reactiontime="0" swimtime="00:06:34.76" resultid="5350" heatid="4949" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.24" />
                    <SPLIT distance="100" swimtime="00:01:40.57" />
                    <SPLIT distance="150" swimtime="00:02:32.19" />
                    <SPLIT distance="200" swimtime="00:03:24.56" />
                    <SPLIT distance="250" swimtime="00:04:17.69" />
                    <SPLIT distance="300" swimtime="00:05:08.50" />
                    <SPLIT distance="350" swimtime="00:05:52.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaella" lastname="Guerra" birthdate="2012-04-02" gender="F" nation="BRA" license="378337" swrid="5603850" athleteid="4617" externalid="378337">
              <RESULTS>
                <RESULT eventid="1093" points="143" reactiontime="0" swimtime="00:00:48.27" resultid="5363" heatid="4862" lane="7" />
                <RESULT eventid="1061" points="136" reactiontime="0" swimtime="00:03:56.79" resultid="5364" heatid="4850" lane="3" />
                <RESULT eventid="1229" points="157" reactiontime="0" swimtime="00:07:13.13" resultid="5365" heatid="4908" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.91" />
                    <SPLIT distance="100" swimtime="00:01:44.43" />
                    <SPLIT distance="150" swimtime="00:02:40.96" />
                    <SPLIT distance="200" swimtime="00:03:36.67" />
                    <SPLIT distance="250" swimtime="00:04:30.04" />
                    <SPLIT distance="300" swimtime="00:05:22.86" />
                    <SPLIT distance="350" swimtime="00:06:19.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1261" points="158" reactiontime="0" swimtime="00:00:42.34" resultid="5366" heatid="4920" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Andre Pangracio" birthdate="2004-01-24" gender="M" nation="BRA" license="265377" swrid="5181504" athleteid="4607" externalid="265377">
              <RESULTS>
                <RESULT eventid="1075" points="440" reactiontime="0" swimtime="00:02:24.05" resultid="5355" heatid="4856" lane="5" entrytime="00:02:16.22" />
                <RESULT eventid="1183" points="434" reactiontime="0" swimtime="00:00:32.95" resultid="5356" heatid="4900" lane="4" entrytime="00:00:30.96" />
                <RESULT eventid="1243" points="459" reactiontime="0" swimtime="00:02:35.73" resultid="5357" heatid="4912" lane="5" entrytime="00:02:26.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="100" swimtime="00:01:13.29" />
                    <SPLIT distance="150" swimtime="00:01:54.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1339" points="453" reactiontime="0" swimtime="00:05:05.63" resultid="5358" heatid="4949" lane="4" entrytime="00:04:51.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                    <SPLIT distance="100" swimtime="00:01:07.55" />
                    <SPLIT distance="150" swimtime="00:01:48.61" />
                    <SPLIT distance="200" swimtime="00:02:28.78" />
                    <SPLIT distance="250" swimtime="00:03:10.69" />
                    <SPLIT distance="300" swimtime="00:03:54.33" />
                    <SPLIT distance="350" swimtime="00:04:30.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Britto" birthdate="2012-10-04" gender="M" nation="BRA" license="378350" swrid="5588566" athleteid="4661" externalid="378350">
              <RESULTS>
                <RESULT eventid="1096" points="138" reactiontime="0" swimtime="00:00:42.91" resultid="5398" heatid="4865" lane="7" entrytime="00:00:51.47" />
                <RESULT eventid="1064" points="147" reactiontime="0" swimtime="00:03:27.54" resultid="5399" heatid="4852" lane="4" entrytime="00:04:42.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.96" />
                    <SPLIT distance="100" swimtime="00:01:37.50" />
                    <SPLIT distance="150" swimtime="00:02:37.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="139" reactiontime="0" swimtime="00:06:49.05" resultid="5400" heatid="4909" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.93" />
                    <SPLIT distance="100" swimtime="00:01:36.64" />
                    <SPLIT distance="150" swimtime="00:02:30.70" />
                    <SPLIT distance="200" swimtime="00:03:23.95" />
                    <SPLIT distance="250" swimtime="00:04:16.16" />
                    <SPLIT distance="300" swimtime="00:05:09.40" />
                    <SPLIT distance="350" swimtime="00:06:02.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="119" reactiontime="0" swimtime="00:00:40.90" resultid="5401" heatid="4925" lane="6" entrytime="00:00:45.05" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Moreschi" birthdate="2012-08-09" gender="M" nation="BRA" license="385715" swrid="5603876" athleteid="4724" externalid="385715">
              <RESULTS>
                <RESULT eventid="1124" points="134" reactiontime="0" swimtime="00:01:27.54" resultid="5448" heatid="4878" lane="6" entrytime="00:01:46.68" />
                <RESULT eventid="1172" points="116" reactiontime="0" swimtime="00:00:51.06" resultid="5449" heatid="4896" lane="2" entrytime="00:00:59.00" />
                <RESULT eventid="1232" points="138" reactiontime="0" swimtime="00:06:49.79" resultid="5450" heatid="4909" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.84" />
                    <SPLIT distance="100" swimtime="00:01:36.79" />
                    <SPLIT distance="150" swimtime="00:02:30.80" />
                    <SPLIT distance="200" swimtime="00:03:25.20" />
                    <SPLIT distance="250" swimtime="00:04:16.89" />
                    <SPLIT distance="300" swimtime="00:05:10.32" />
                    <SPLIT distance="350" swimtime="00:06:03.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="111" reactiontime="0" swimtime="00:01:54.76" resultid="5451" heatid="4953" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mirella" lastname="Paula Correia Thomé" birthdate="2012-02-12" gender="F" nation="BRA" license="382236" swrid="5603886" athleteid="4700" externalid="382236">
              <RESULTS>
                <RESULT eventid="1093" points="133" reactiontime="0" swimtime="00:00:49.45" resultid="5429" heatid="4862" lane="3" entrytime="00:00:52.41" />
                <RESULT eventid="1061" points="70" reactiontime="0" swimtime="00:04:55.20" resultid="5430" heatid="4851" lane="7" />
                <RESULT eventid="1229" points="160" reactiontime="0" swimtime="00:07:10.39" resultid="5431" heatid="4908" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.62" />
                    <SPLIT distance="100" swimtime="00:01:41.50" />
                    <SPLIT distance="150" swimtime="00:02:37.78" />
                    <SPLIT distance="200" swimtime="00:03:32.00" />
                    <SPLIT distance="250" swimtime="00:04:30.31" />
                    <SPLIT distance="300" swimtime="00:05:20.82" />
                    <SPLIT distance="350" swimtime="00:06:16.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1309" points="101" reactiontime="0" swimtime="00:00:52.29" resultid="5432" heatid="4940" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benicio" lastname="Garcia" birthdate="2011-09-09" gender="M" nation="BRA" license="378347" swrid="5603842" athleteid="4651" externalid="378347">
              <RESULTS>
                <RESULT eventid="1096" points="176" reactiontime="0" swimtime="00:00:39.60" resultid="5390" heatid="4865" lane="5" entrytime="00:00:43.13" />
                <RESULT eventid="1124" points="170" reactiontime="0" swimtime="00:01:20.91" resultid="5391" heatid="4879" lane="6" entrytime="00:01:23.84" />
                <RESULT eventid="1232" points="182" reactiontime="0" swimtime="00:06:14.24" resultid="5392" heatid="4909" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.36" />
                    <SPLIT distance="100" swimtime="00:01:28.91" />
                    <SPLIT distance="150" swimtime="00:02:17.64" />
                    <SPLIT distance="200" swimtime="00:03:04.95" />
                    <SPLIT distance="250" swimtime="00:03:53.15" />
                    <SPLIT distance="300" swimtime="00:04:41.05" />
                    <SPLIT distance="350" swimtime="00:05:29.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="176" reactiontime="0" swimtime="00:00:35.93" resultid="5393" heatid="4925" lane="4" entrytime="00:00:40.12" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Magalhães Rezende" birthdate="2010-05-29" gender="F" nation="BRA" license="366960" swrid="5588793" athleteid="4592" externalid="366960">
              <RESULTS>
                <RESULT eventid="1067" points="342" reactiontime="0" swimtime="00:02:54.23" resultid="5343" heatid="4853" lane="5" entrytime="00:03:15.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                    <SPLIT distance="100" swimtime="00:01:23.62" />
                    <SPLIT distance="150" swimtime="00:02:15.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="348" reactiontime="0" swimtime="00:11:21.08" resultid="5344" heatid="4901" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:11:22.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1235" points="321" reactiontime="0" swimtime="00:03:16.51" resultid="5345" heatid="4910" lane="4" />
                <RESULT eventid="1315" points="312" reactiontime="0" swimtime="00:00:35.94" resultid="5346" heatid="4944" lane="2" entrytime="00:00:37.47" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Rezende" birthdate="2012-01-23" gender="F" nation="BRA" license="370669" swrid="5603899" athleteid="4690" externalid="370669">
              <RESULTS>
                <RESULT eventid="1061" points="163" reactiontime="0" swimtime="00:03:43.07" resultid="5421" heatid="4851" lane="3" entrytime="00:04:02.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.78" />
                    <SPLIT distance="100" swimtime="00:01:51.89" />
                    <SPLIT distance="150" swimtime="00:02:52.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1169" points="182" reactiontime="0" swimtime="00:00:50.35" resultid="5422" heatid="4894" lane="3" entrytime="00:00:51.84" />
                <RESULT eventid="1261" points="208" reactiontime="0" swimtime="00:00:38.69" resultid="5423" heatid="4922" lane="2" entrytime="00:00:44.73" />
                <RESULT eventid="1347" points="165" reactiontime="0" swimtime="00:01:53.50" resultid="5424" heatid="4951" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theodoro" lastname="Marques Serra" birthdate="2009-11-24" gender="M" nation="BRA" license="370661" swrid="5603870" athleteid="4685" externalid="370661">
              <RESULTS>
                <RESULT eventid="1075" reactiontime="0" status="DSQ" swimtime="00:00:00.00" resultid="5417" heatid="4854" lane="3" />
                <RESULT eventid="1107" points="206" reactiontime="0" swimtime="00:00:37.61" resultid="5418" heatid="4868" lane="3" entrytime="00:00:39.23" />
                <RESULT eventid="1275" points="261" reactiontime="0" swimtime="00:00:31.51" resultid="5419" heatid="4931" lane="6" entrytime="00:00:31.90" />
                <RESULT eventid="1291" points="233" reactiontime="0" swimtime="00:02:51.50" resultid="5420" heatid="4934" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.12" />
                    <SPLIT distance="100" swimtime="00:01:22.47" />
                    <SPLIT distance="150" swimtime="00:02:07.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Rossi" birthdate="2012-05-21" gender="M" nation="BRA" license="378346" swrid="5603901" athleteid="4646" externalid="378346">
              <RESULTS>
                <RESULT eventid="1096" points="94" reactiontime="0" swimtime="00:00:48.70" resultid="5386" heatid="4863" lane="4" />
                <RESULT eventid="1124" points="154" reactiontime="0" swimtime="00:01:23.57" resultid="5387" heatid="4878" lane="7" entrytime="00:02:00.51" />
                <RESULT eventid="1264" points="150" reactiontime="0" swimtime="00:00:37.91" resultid="5388" heatid="4925" lane="7" entrytime="00:00:51.08" />
                <RESULT eventid="1312" points="111" reactiontime="0" swimtime="00:00:45.18" resultid="5389" heatid="4942" lane="5" entrytime="00:01:10.59" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15981" nation="BRA" clubid="4142" swrid="93783" name="Quinto Nado" shortname="5º Nado">
          <ATHLETES>
            <ATHLETE firstname="Gabriela" lastname="Gomes" birthdate="2011-12-03" gender="F" nation="BRA" license="382051" swrid="5603846" athleteid="4184" externalid="382051">
              <RESULTS>
                <RESULT eventid="1389" points="135" reactiontime="0" swimtime="00:01:46.81" resultid="5013" heatid="4961" lane="5" entrytime="00:02:08.74" />
                <RESULT eventid="1417" points="158" reactiontime="0" swimtime="00:03:23.95" resultid="5014" heatid="4967" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.20" />
                    <SPLIT distance="100" swimtime="00:01:41.01" />
                    <SPLIT distance="150" swimtime="00:02:33.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Takemura Couto" birthdate="2010-02-08" gender="F" nation="BRA" license="376950" swrid="5603919" athleteid="4171" externalid="376950">
              <RESULTS>
                <RESULT eventid="1067" points="279" reactiontime="0" swimtime="00:03:06.28" resultid="5002" heatid="4853" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.24" />
                    <SPLIT distance="100" swimtime="00:01:26.03" />
                    <SPLIT distance="150" swimtime="00:02:22.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="321" reactiontime="0" swimtime="00:01:13.38" resultid="5003" heatid="4880" lane="5" entrytime="00:01:14.23" />
                <RESULT eventid="1213" points="289" reactiontime="0" swimtime="00:05:53.71" resultid="5004" heatid="4906" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:05:55.57" />
                    <SPLIT distance="100" swimtime="00:06:03.81" />
                    <SPLIT distance="150" swimtime="00:06:12.45" />
                    <SPLIT distance="200" swimtime="00:06:12.65" />
                    <SPLIT distance="250" swimtime="00:06:12.87" />
                    <SPLIT distance="300" swimtime="00:06:13.08" />
                    <SPLIT distance="350" swimtime="00:06:13.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1283" reactiontime="0" status="DSQ" swimtime="00:00:00.00" resultid="5005" heatid="4933" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.41" />
                    <SPLIT distance="100" swimtime="00:01:26.32" />
                    <SPLIT distance="150" swimtime="00:02:12.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1353" points="292" reactiontime="0" swimtime="00:02:46.20" resultid="5006" heatid="4954" lane="3" entrytime="00:03:00.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.46" />
                    <SPLIT distance="100" swimtime="00:01:20.20" />
                    <SPLIT distance="150" swimtime="00:02:05.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1395" points="293" reactiontime="0" swimtime="00:01:22.64" resultid="5007" heatid="4963" lane="3" entrytime="00:01:24.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Vieira Daudt" birthdate="2014-09-29" gender="M" nation="BRA" license="392039" swrid="5603927" athleteid="4198" externalid="392039">
              <RESULTS>
                <RESULT eventid="1166" points="41" reactiontime="0" swimtime="00:01:11.78" resultid="5024" heatid="4891" lane="5" />
                <RESULT eventid="1258" points="59" reactiontime="0" swimtime="00:00:51.57" resultid="5025" heatid="4919" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Betina" lastname="Queiroz" birthdate="2007-09-11" gender="F" nation="BRA" license="357155" swrid="5603897" athleteid="4157" externalid="357155">
              <RESULTS>
                <RESULT eventid="1127" points="505" reactiontime="0" swimtime="00:01:03.09" resultid="4990" heatid="4881" lane="5" entrytime="00:01:03.85" />
                <RESULT eventid="1191" points="476" reactiontime="0" swimtime="00:10:13.83" resultid="4991" heatid="4901" lane="4" entrytime="00:10:16.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:10:20.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="487" reactiontime="0" swimtime="00:04:57.16" resultid="4992" heatid="4906" lane="4" entrytime="00:04:52.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                    <SPLIT distance="100" swimtime="00:01:10.43" />
                    <SPLIT distance="150" swimtime="00:01:47.60" />
                    <SPLIT distance="200" swimtime="00:02:25.62" />
                    <SPLIT distance="250" swimtime="00:03:04.08" />
                    <SPLIT distance="300" swimtime="00:03:42.30" />
                    <SPLIT distance="350" swimtime="00:04:20.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="423" reactiontime="0" swimtime="00:00:30.53" resultid="4993" heatid="4928" lane="3" entrytime="00:00:30.34" />
                <RESULT eventid="1353" points="475" reactiontime="0" swimtime="00:02:21.34" resultid="4994" heatid="4955" lane="4" entrytime="00:02:18.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                    <SPLIT distance="100" swimtime="00:01:08.03" />
                    <SPLIT distance="150" swimtime="00:01:44.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1445" points="301" reactiontime="0" swimtime="00:01:21.39" resultid="4995" heatid="4974" lane="6" entrytime="00:01:28.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco" lastname="Silva Telles" birthdate="2011-07-19" gender="M" nation="BRA" license="377311" swrid="5603911" athleteid="4178" externalid="377311">
              <RESULTS>
                <RESULT eventid="1124" points="134" reactiontime="0" swimtime="00:01:27.57" resultid="5008" heatid="4878" lane="5" entrytime="00:01:40.10" />
                <RESULT eventid="1172" reactiontime="0" status="DSQ" swimtime="00:00:00.00" resultid="5009" heatid="4896" lane="6" entrytime="00:00:52.56" />
                <RESULT eventid="1264" points="137" reactiontime="0" swimtime="00:00:39.08" resultid="5010" heatid="4925" lane="3" entrytime="00:00:43.18" />
                <RESULT eventid="1350" points="126" reactiontime="0" swimtime="00:01:50.09" resultid="5011" heatid="4953" lane="3" entrytime="00:02:02.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1420" points="123" reactiontime="0" swimtime="00:03:19.61" resultid="5012" heatid="4968" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.09" />
                    <SPLIT distance="100" swimtime="00:01:32.63" />
                    <SPLIT distance="150" swimtime="00:02:27.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Clara Bobroff" birthdate="2013-02-09" gender="F" nation="BRA" license="391752" swrid="5419807" athleteid="4194" externalid="391752">
              <RESULTS>
                <RESULT eventid="1115" points="156" reactiontime="0" swimtime="00:01:33.29" resultid="5021" heatid="4870" lane="5" />
                <RESULT eventid="1163" points="133" reactiontime="0" swimtime="00:00:55.85" resultid="5022" heatid="4889" lane="3" />
                <RESULT eventid="1255" points="167" reactiontime="0" swimtime="00:00:41.58" resultid="5023" heatid="4914" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Bordini Zocco" birthdate="2008-08-04" gender="F" nation="BRA" license="385677" swrid="5332871" athleteid="4187" externalid="385677">
              <RESULTS>
                <RESULT eventid="1067" points="295" reactiontime="0" swimtime="00:03:02.87" resultid="5015" heatid="4853" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.19" />
                    <SPLIT distance="100" swimtime="00:01:26.39" />
                    <SPLIT distance="150" swimtime="00:02:21.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="331" reactiontime="0" swimtime="00:01:12.57" resultid="5016" heatid="4880" lane="6" entrytime="00:01:18.54" />
                <RESULT eventid="1213" points="328" reactiontime="0" swimtime="00:05:38.99" resultid="5017" heatid="4906" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.96" />
                    <SPLIT distance="100" swimtime="00:01:20.54" />
                    <SPLIT distance="150" swimtime="00:02:03.75" />
                    <SPLIT distance="200" swimtime="00:02:47.75" />
                    <SPLIT distance="250" swimtime="00:03:31.10" />
                    <SPLIT distance="300" swimtime="00:04:15.16" />
                    <SPLIT distance="350" swimtime="00:04:59.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="305" reactiontime="0" swimtime="00:00:34.04" resultid="5018" heatid="4927" lane="5" entrytime="00:00:34.98" />
                <RESULT eventid="1369" points="265" reactiontime="0" swimtime="00:01:37.03" resultid="5019" heatid="4958" lane="5" entrytime="00:01:46.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="298" reactiontime="0" swimtime="00:01:24.52" resultid="5020" heatid="4970" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Poletti Veiga" birthdate="2010-10-01" gender="F" nation="BRA" license="376951" swrid="5603895" athleteid="4150" externalid="376951">
              <RESULTS>
                <RESULT eventid="1067" reactiontime="0" status="DSQ" swimtime="00:00:00.00" resultid="4984" heatid="4853" lane="6" />
                <RESULT eventid="1127" points="353" reactiontime="0" swimtime="00:01:11.06" resultid="4985" heatid="4880" lane="3" entrytime="00:01:17.92" />
                <RESULT eventid="1213" points="370" reactiontime="0" swimtime="00:05:25.59" resultid="4986" heatid="4906" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.62" />
                    <SPLIT distance="100" swimtime="00:01:17.84" />
                    <SPLIT distance="150" swimtime="00:01:59.02" />
                    <SPLIT distance="200" swimtime="00:02:41.36" />
                    <SPLIT distance="250" swimtime="00:03:23.54" />
                    <SPLIT distance="300" swimtime="00:04:04.89" />
                    <SPLIT distance="350" swimtime="00:04:47.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="364" reactiontime="0" swimtime="00:00:32.09" resultid="4987" heatid="4927" lane="4" entrytime="00:00:34.46" />
                <RESULT eventid="1353" points="361" reactiontime="0" swimtime="00:02:34.79" resultid="4988" heatid="4954" lane="5" entrytime="00:02:54.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.86" />
                    <SPLIT distance="100" swimtime="00:01:15.49" />
                    <SPLIT distance="150" swimtime="00:01:56.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1395" points="293" reactiontime="0" swimtime="00:01:22.59" resultid="4989" heatid="4963" lane="6" entrytime="00:01:31.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Kikuchi Fujii" birthdate="2007-01-04" gender="M" nation="BRA" license="297805" swrid="5603863" athleteid="4143" externalid="297805">
              <RESULTS>
                <RESULT eventid="1075" reactiontime="0" status="DSQ" swimtime="00:00:00.00" resultid="4978" heatid="4856" lane="3" entrytime="00:02:16.93" />
                <RESULT eventid="1183" points="508" reactiontime="0" swimtime="00:00:31.25" resultid="4979" heatid="4900" lane="3" entrytime="00:00:33.52" />
                <RESULT eventid="1243" reactiontime="0" status="DSQ" swimtime="00:00:00.00" resultid="4980" heatid="4912" lane="3" entrytime="00:02:26.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="100" swimtime="00:01:08.99" />
                    <SPLIT distance="150" swimtime="00:01:46.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1323" points="495" reactiontime="0" swimtime="00:00:27.49" resultid="4981" heatid="4945" lane="3" />
                <RESULT eventid="1377" points="587" reactiontime="0" swimtime="00:01:05.99" resultid="4982" heatid="4960" lane="4" entrytime="00:01:07.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="451" reactiontime="0" swimtime="00:01:02.26" resultid="4983" heatid="4976" lane="5" entrytime="00:01:02.31" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Vieira Daudt" birthdate="2008-08-14" gender="M" nation="BRA" license="350467" swrid="5603926" athleteid="4164" externalid="350467">
              <RESULTS>
                <RESULT eventid="1075" points="263" reactiontime="0" swimtime="00:02:51.08" resultid="4996" heatid="4855" lane="2" />
                <RESULT eventid="1135" points="312" reactiontime="0" swimtime="00:01:06.05" resultid="4997" heatid="4884" lane="7" entrytime="00:01:09.11" />
                <RESULT eventid="1221" points="281" reactiontime="0" swimtime="00:05:23.89" resultid="4998" heatid="4907" lane="5" entrytime="00:05:53.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.79" />
                    <SPLIT distance="100" swimtime="00:01:18.86" />
                    <SPLIT distance="150" swimtime="00:01:58.82" />
                    <SPLIT distance="200" swimtime="00:02:40.21" />
                    <SPLIT distance="250" swimtime="00:03:20.08" />
                    <SPLIT distance="300" swimtime="00:04:02.23" />
                    <SPLIT distance="350" swimtime="00:04:42.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1291" points="264" reactiontime="0" swimtime="00:02:44.59" resultid="4999" heatid="4934" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                    <SPLIT distance="100" swimtime="00:01:21.21" />
                    <SPLIT distance="150" swimtime="00:02:03.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1403" points="271" reactiontime="0" swimtime="00:01:14.61" resultid="5000" heatid="4964" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="220" reactiontime="0" swimtime="00:01:19.11" resultid="5001" heatid="4975" lane="5" entrytime="00:01:33.68" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2416" nation="BRA" clubid="4201" swrid="93758" name="Associação de Pais e Atletas de Natação de Maringá" shortname="Apan/Maringá">
          <ATHLETES>
            <ATHLETE firstname="Julia" lastname="Vitoria Moreira Ferreira" birthdate="2012-08-04" gender="F" nation="BRA" license="392098" swrid="5603928" athleteid="4496" externalid="392098">
              <RESULTS>
                <RESULT eventid="1093" reactiontime="0" status="DSQ" swimtime="00:00:00.00" resultid="5267" heatid="4861" lane="4" />
                <RESULT eventid="1169" points="39" reactiontime="0" swimtime="00:01:23.55" resultid="5268" heatid="4893" lane="5" />
                <RESULT eventid="1261" points="43" reactiontime="0" swimtime="00:01:05.44" resultid="5269" heatid="4921" lane="2" />
                <RESULT eventid="1347" points="44" reactiontime="0" swimtime="00:02:55.59" resultid="5270" heatid="4950" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Muniz" birthdate="2012-09-03" gender="M" nation="BRA" license="392106" swrid="5603877" athleteid="4533" externalid="392106">
              <RESULTS>
                <RESULT eventid="1124" points="30" reactiontime="0" swimtime="00:02:23.27" resultid="5296" heatid="4877" lane="2" />
                <RESULT eventid="1172" points="23" reactiontime="0" swimtime="00:01:26.78" resultid="5297" heatid="4895" lane="3" />
                <RESULT eventid="1264" points="36" reactiontime="0" swimtime="00:01:00.66" resultid="5298" heatid="4923" lane="2" />
                <RESULT eventid="1350" points="27" reactiontime="0" swimtime="00:03:03.11" resultid="5299" heatid="4952" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Stephany" birthdate="2012-07-27" gender="F" nation="BRA" license="382210" swrid="5603917" athleteid="4434" externalid="382210">
              <RESULTS>
                <RESULT eventid="1093" points="123" reactiontime="0" swimtime="00:00:50.69" resultid="5216" heatid="4862" lane="6" entrytime="00:01:00.33" />
                <RESULT eventid="1121" points="137" reactiontime="0" swimtime="00:01:37.45" resultid="5217" heatid="4875" lane="2" entrytime="00:01:54.49" />
                <RESULT eventid="1261" points="164" reactiontime="0" swimtime="00:00:41.82" resultid="5218" heatid="4921" lane="5" entrytime="00:00:52.31" />
                <RESULT eventid="1309" points="97" reactiontime="0" swimtime="00:00:52.90" resultid="5219" heatid="4941" lane="3" entrytime="00:01:02.99" />
                <RESULT eventid="1417" points="129" reactiontime="0" swimtime="00:03:37.88" resultid="5220" heatid="4967" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.90" />
                    <SPLIT distance="100" swimtime="00:01:44.17" />
                    <SPLIT distance="150" swimtime="00:02:41.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" reactiontime="0" status="DSQ" swimtime="00:00:00.00" resultid="5221" heatid="4972" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juan" lastname="Bernardo Padua" birthdate="2013-07-15" gender="M" nation="BRA" license="392108" swrid="5305422" athleteid="4543" externalid="392108">
              <RESULTS>
                <RESULT eventid="1118" points="50" reactiontime="0" swimtime="00:02:01.04" resultid="5304" heatid="4872" lane="3" />
                <RESULT eventid="1166" points="50" reactiontime="0" swimtime="00:01:07.45" resultid="5305" heatid="4892" lane="6" />
                <RESULT eventid="1258" points="56" reactiontime="0" swimtime="00:00:52.65" resultid="5306" heatid="4919" lane="2" />
                <RESULT eventid="1306" points="27" reactiontime="0" swimtime="00:01:12.47" resultid="5307" heatid="4938" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Pacheco" birthdate="2006-12-20" gender="M" nation="BRA" license="336850" swrid="5603854" athleteid="4259" externalid="336850">
              <RESULTS>
                <RESULT eventid="1075" points="403" reactiontime="0" swimtime="00:02:28.41" resultid="5070" heatid="4856" lane="6" entrytime="00:02:29.55" />
                <RESULT eventid="1151" points="294" reactiontime="0" swimtime="00:02:42.78" resultid="5071" heatid="4887" lane="4" entrytime="00:02:34.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                    <SPLIT distance="100" swimtime="00:01:14.88" />
                    <SPLIT distance="150" swimtime="00:01:57.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1339" points="393" reactiontime="0" swimtime="00:05:20.37" resultid="5072" heatid="4949" lane="5" entrytime="00:05:28.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                    <SPLIT distance="100" swimtime="00:01:10.42" />
                    <SPLIT distance="150" swimtime="00:01:52.99" />
                    <SPLIT distance="200" swimtime="00:02:34.63" />
                    <SPLIT distance="250" swimtime="00:03:22.59" />
                    <SPLIT distance="300" swimtime="00:04:09.83" />
                    <SPLIT distance="350" swimtime="00:04:46.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="405" reactiontime="0" swimtime="00:01:04.56" resultid="5073" heatid="4976" lane="3" entrytime="00:01:05.62" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Oliveira Silva" birthdate="2013-02-05" gender="M" nation="BRA" license="392109" swrid="5603880" athleteid="4548" externalid="392109" />
            <ATHLETE firstname="Matheus" lastname="Gongora De Campos" birthdate="2013-02-17" gender="M" nation="BRA" license="377262" swrid="5603847" athleteid="4390" externalid="377262">
              <RESULTS>
                <RESULT eventid="1090" points="127" reactiontime="0" swimtime="00:00:44.18" resultid="5179" heatid="4860" lane="4" entrytime="00:00:45.23" />
                <RESULT eventid="1118" points="128" reactiontime="0" swimtime="00:01:28.76" resultid="5180" heatid="4873" lane="4" entrytime="00:01:31.49" />
                <RESULT eventid="1210" points="105" reactiontime="0" swimtime="00:01:44.27" resultid="5181" heatid="4905" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="119" reactiontime="0" swimtime="00:00:40.91" resultid="5182" heatid="4919" lane="4" entrytime="00:00:42.61" />
                <RESULT eventid="1414" points="139" reactiontime="0" swimtime="00:03:11.74" resultid="5183" heatid="4966" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.82" />
                    <SPLIT distance="100" swimtime="00:01:37.05" />
                    <SPLIT distance="150" swimtime="00:02:25.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wellington" lastname="De Lima" birthdate="2008-03-01" gender="M" nation="BRA" license="370024" swrid="5470912" athleteid="4215" externalid="370024">
              <RESULTS>
                <RESULT eventid="1135" points="443" reactiontime="0" swimtime="00:00:58.80" resultid="5036" heatid="4884" lane="4" entrytime="00:00:59.80" />
                <RESULT eventid="1275" points="379" reactiontime="0" swimtime="00:00:27.84" resultid="5037" heatid="4932" lane="6" entrytime="00:00:27.67" />
                <RESULT eventid="1323" points="290" reactiontime="0" swimtime="00:00:32.84" resultid="5038" heatid="4945" lane="5" />
                <RESULT eventid="1361" points="376" reactiontime="0" swimtime="00:02:17.56" resultid="5039" heatid="4957" lane="6" entrytime="00:02:17.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                    <SPLIT distance="100" swimtime="00:01:05.33" />
                    <SPLIT distance="150" swimtime="00:01:41.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1403" points="258" reactiontime="0" swimtime="00:01:15.89" resultid="5040" heatid="4964" lane="4" entrytime="00:01:14.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Pavão" birthdate="2012-04-04" gender="F" nation="BRA" license="377259" swrid="5603888" athleteid="4371" externalid="377259">
              <RESULTS>
                <RESULT eventid="1093" points="158" reactiontime="0" swimtime="00:00:46.71" resultid="5163" heatid="4862" lane="4" entrytime="00:00:48.08" />
                <RESULT eventid="1061" points="151" reactiontime="0" swimtime="00:03:48.66" resultid="5164" heatid="4851" lane="2" entrytime="00:04:11.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.77" />
                    <SPLIT distance="100" swimtime="00:01:52.61" />
                    <SPLIT distance="150" swimtime="00:02:54.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1261" points="159" reactiontime="0" swimtime="00:00:42.29" resultid="5165" heatid="4922" lane="7" entrytime="00:00:45.69" />
                <RESULT eventid="1389" reactiontime="0" status="DSQ" swimtime="00:00:00.00" resultid="5166" heatid="4961" lane="3" />
                <RESULT eventid="1417" points="127" reactiontime="0" swimtime="00:03:39.26" resultid="5167" heatid="4967" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.46" />
                    <SPLIT distance="100" swimtime="00:01:45.36" />
                    <SPLIT distance="150" swimtime="00:02:44.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Diego" lastname="Duarte Rezende" birthdate="2006-01-25" gender="M" nation="BRA" license="313013" swrid="5498173" athleteid="4246" externalid="313013">
              <RESULTS>
                <RESULT eventid="1107" points="438" reactiontime="0" swimtime="00:00:29.25" resultid="5060" heatid="4868" lane="4" entrytime="00:00:28.97" />
                <RESULT eventid="1135" points="490" reactiontime="0" swimtime="00:00:56.86" resultid="5061" heatid="4885" lane="2" entrytime="00:00:57.85" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabrielle" lastname="Borba" birthdate="2014-06-15" gender="F" nation="BRA" license="385705" swrid="5323267" athleteid="4447" externalid="385705">
              <RESULTS>
                <RESULT eventid="1087" points="76" reactiontime="0" swimtime="00:00:59.60" resultid="5227" heatid="4858" lane="5" />
                <RESULT eventid="1163" points="72" reactiontime="0" swimtime="00:01:08.61" resultid="5228" heatid="4889" lane="4" />
                <RESULT eventid="1255" points="97" reactiontime="0" swimtime="00:00:49.81" resultid="5229" heatid="4915" lane="5" />
                <RESULT eventid="1303" points="71" reactiontime="0" swimtime="00:00:58.61" resultid="5230" heatid="4936" lane="4" />
                <RESULT eventid="1411" points="93" reactiontime="0" swimtime="00:04:03.21" resultid="5231" heatid="4965" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.58" />
                    <SPLIT distance="100" swimtime="00:01:57.60" />
                    <SPLIT distance="150" swimtime="00:03:01.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Donato De Morais" birthdate="2009-03-28" gender="F" nation="BRA" license="345588" swrid="5485198" athleteid="4274" externalid="345588">
              <RESULTS>
                <RESULT eventid="1099" points="346" reactiontime="0" swimtime="00:00:35.98" resultid="5082" heatid="4866" lane="5" entrytime="00:00:37.33" />
                <RESULT eventid="1191" points="345" reactiontime="0" swimtime="00:11:23.15" resultid="5083" heatid="4901" lane="5" entrytime="00:10:59.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:11:24.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1283" points="354" reactiontime="0" swimtime="00:02:48.05" resultid="5084" heatid="4933" lane="5" entrytime="00:02:44.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                    <SPLIT distance="100" swimtime="00:01:22.31" />
                    <SPLIT distance="150" swimtime="00:02:06.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1395" points="346" reactiontime="0" swimtime="00:01:18.15" resultid="5085" heatid="4963" lane="4" entrytime="00:01:16.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1423" points="290" reactiontime="0" swimtime="00:01:25.35" resultid="5086" heatid="4970" lane="4" entrytime="00:01:58.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lavinia" lastname="Bossoni" birthdate="2013-11-03" gender="F" nation="BRA" license="377260" swrid="5343093" athleteid="4377" externalid="377260">
              <RESULTS>
                <RESULT eventid="1087" points="152" reactiontime="0" swimtime="00:00:47.25" resultid="5168" heatid="4859" lane="3" entrytime="00:00:54.12" />
                <RESULT eventid="1163" points="122" reactiontime="0" swimtime="00:00:57.54" resultid="5169" heatid="4890" lane="5" entrytime="00:01:03.15" />
                <RESULT eventid="1207" points="151" reactiontime="0" swimtime="00:01:46.09" resultid="5170" heatid="4904" lane="3" />
                <RESULT eventid="1255" points="136" reactiontime="0" swimtime="00:00:44.54" resultid="5171" heatid="4916" lane="3" entrytime="00:00:48.51" />
                <RESULT eventid="1411" points="114" reactiontime="0" swimtime="00:03:46.94" resultid="5172" heatid="4965" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.52" />
                    <SPLIT distance="100" swimtime="00:01:50.00" />
                    <SPLIT distance="150" swimtime="00:02:50.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="José Da Silva" birthdate="2008-04-04" gender="M" nation="BRA" license="318192" swrid="5603858" athleteid="4209" externalid="318192">
              <RESULTS>
                <RESULT eventid="1135" points="572" reactiontime="0" swimtime="00:00:54.00" resultid="5031" heatid="4885" lane="3" entrytime="00:00:55.23" />
                <RESULT eventid="1221" points="488" reactiontime="0" swimtime="00:04:29.42" resultid="5032" heatid="4907" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                    <SPLIT distance="100" swimtime="00:01:06.01" />
                    <SPLIT distance="150" swimtime="00:01:40.24" />
                    <SPLIT distance="200" swimtime="00:02:14.84" />
                    <SPLIT distance="250" swimtime="00:02:49.64" />
                    <SPLIT distance="300" swimtime="00:03:23.83" />
                    <SPLIT distance="350" swimtime="00:03:58.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1275" points="525" reactiontime="0" swimtime="00:00:24.98" resultid="5033" heatid="4932" lane="5" entrytime="00:00:25.18" />
                <RESULT eventid="1361" points="582" reactiontime="0" swimtime="00:01:59.00" resultid="5034" heatid="4957" lane="5" entrytime="00:02:07.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.21" />
                    <SPLIT distance="100" swimtime="00:00:57.16" />
                    <SPLIT distance="150" swimtime="00:01:27.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="519" reactiontime="0" swimtime="00:00:59.45" resultid="5035" heatid="4976" lane="4" entrytime="00:01:00.24" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Santos Carraro" birthdate="2014-06-04" gender="M" nation="BRA" license="392097" swrid="5603908" athleteid="4490" externalid="392097">
              <RESULTS>
                <RESULT eventid="1090" points="67" reactiontime="0" swimtime="00:00:54.44" resultid="5262" heatid="4860" lane="6" />
                <RESULT eventid="1118" points="77" reactiontime="0" swimtime="00:01:45.24" resultid="5263" heatid="4872" lane="5" />
                <RESULT eventid="1258" points="81" reactiontime="0" swimtime="00:00:46.53" resultid="5264" heatid="4918" lane="3" />
                <RESULT eventid="1306" points="54" reactiontime="0" swimtime="00:00:57.46" resultid="5265" heatid="4939" lane="4" />
                <RESULT eventid="1414" points="75" reactiontime="0" swimtime="00:03:55.23" resultid="5266" heatid="4966" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.48" />
                    <SPLIT distance="100" swimtime="00:01:51.55" />
                    <SPLIT distance="150" swimtime="00:02:56.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Campelo" birthdate="2011-09-12" gender="M" nation="BRA" license="366963" swrid="5588742" athleteid="4322" externalid="366963">
              <RESULTS>
                <RESULT eventid="1096" reactiontime="0" status="DNS" swimtime="00:00:00.00" resultid="5122" entrytime="00:00:38.81" />
                <RESULT eventid="1124" reactiontime="0" status="DNS" swimtime="00:00:00.00" resultid="5123" entrytime="00:01:15.31" />
                <RESULT eventid="1264" reactiontime="0" status="DNS" swimtime="00:00:00.00" resultid="5124" entrytime="00:00:31.26" />
                <RESULT eventid="1312" reactiontime="0" status="DNS" swimtime="00:00:00.00" resultid="5125" entrytime="00:00:35.74" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Schuch Pimpao" birthdate="2010-12-31" gender="M" nation="BRA" license="355586" swrid="5588908" athleteid="4317" externalid="355586">
              <RESULTS>
                <RESULT eventid="1135" points="228" reactiontime="0" swimtime="00:01:13.30" resultid="5118" heatid="4883" lane="3" entrytime="00:01:15.70" />
                <RESULT eventid="1183" points="173" reactiontime="0" swimtime="00:00:44.77" resultid="5119" heatid="4899" lane="5" entrytime="00:00:45.18" />
                <RESULT eventid="1275" points="229" reactiontime="0" swimtime="00:00:32.92" resultid="5120" heatid="4931" lane="2" entrytime="00:00:32.47" />
                <RESULT eventid="1403" points="197" reactiontime="0" swimtime="00:01:23.00" resultid="5121" heatid="4964" lane="3" entrytime="00:01:22.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Forti Francisco" birthdate="2015-07-08" gender="M" nation="BRA" license="392104" swrid="5534395" athleteid="4523" externalid="392104">
              <RESULTS>
                <RESULT eventid="1085" points="32" reactiontime="0" swimtime="00:00:32.44" resultid="5288" heatid="4857" lane="5" />
                <RESULT eventid="1161" points="27" reactiontime="0" swimtime="00:00:38.16" resultid="5289" heatid="4888" lane="5" />
                <RESULT eventid="1253" points="37" reactiontime="0" swimtime="00:00:27.23" resultid="5290" heatid="4913" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Peroni Passafaro" birthdate="2013-09-17" gender="F" nation="BRA" license="370659" swrid="5603893" athleteid="4345" externalid="370659">
              <RESULTS>
                <RESULT eventid="1087" points="140" reactiontime="0" swimtime="00:00:48.65" resultid="5141" heatid="4859" lane="5" entrytime="00:00:51.32" />
                <RESULT eventid="1115" points="123" reactiontime="0" swimtime="00:01:40.99" resultid="5142" heatid="4871" lane="5" entrytime="00:01:44.13" />
                <RESULT eventid="1207" points="129" reactiontime="0" swimtime="00:01:51.72" resultid="5143" heatid="4904" lane="4" entrytime="00:02:29.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1255" points="133" reactiontime="0" swimtime="00:00:44.87" resultid="5144" heatid="4916" lane="4" entrytime="00:00:37.63" />
                <RESULT eventid="1411" points="125" reactiontime="0" swimtime="00:03:40.50" resultid="5145" heatid="4965" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.85" />
                    <SPLIT distance="100" swimtime="00:01:51.01" />
                    <SPLIT distance="150" swimtime="00:02:49.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amanda" lastname="Beatriz Meira" birthdate="2012-04-11" gender="F" nation="BRA" license="392094" swrid="5305414" athleteid="4476" externalid="392094">
              <RESULTS>
                <RESULT eventid="1093" points="46" reactiontime="0" swimtime="00:01:10.45" resultid="5251" heatid="4861" lane="2" />
                <RESULT eventid="1121" points="58" reactiontime="0" swimtime="00:02:09.10" resultid="5252" heatid="4874" lane="4" />
                <RESULT eventid="1261" points="71" reactiontime="0" swimtime="00:00:55.14" resultid="5253" heatid="4921" lane="6" />
                <RESULT eventid="1309" points="42" reactiontime="0" swimtime="00:01:09.74" resultid="5254" heatid="4941" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Biason Santana" birthdate="2009-01-21" gender="M" nation="BRA" license="366969" swrid="5317765" athleteid="4298" externalid="366969">
              <RESULTS>
                <RESULT eventid="1075" points="289" reactiontime="0" swimtime="00:02:45.75" resultid="5102" heatid="4854" lane="4" />
                <RESULT eventid="1135" points="360" reactiontime="0" swimtime="00:01:03.02" resultid="5103" heatid="4884" lane="5" entrytime="00:01:01.56" />
                <RESULT eventid="1275" points="339" reactiontime="0" swimtime="00:00:28.91" resultid="5104" heatid="4932" lane="2" entrytime="00:00:27.71" />
                <RESULT eventid="1323" points="339" reactiontime="0" swimtime="00:00:31.18" resultid="5105" heatid="4947" lane="3" entrytime="00:00:30.69" />
                <RESULT eventid="1361" points="311" reactiontime="0" swimtime="00:02:26.63" resultid="5106" heatid="4957" lane="7" entrytime="00:02:20.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                    <SPLIT distance="100" swimtime="00:01:11.40" />
                    <SPLIT distance="150" swimtime="00:01:48.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="331" reactiontime="0" swimtime="00:01:09.07" resultid="5107" heatid="4976" lane="6" entrytime="00:01:08.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Ayres" birthdate="2012-05-05" gender="M" nation="BRA" license="378035" swrid="5208079" athleteid="4403" externalid="378035">
              <RESULTS>
                <RESULT eventid="1096" points="170" reactiontime="0" swimtime="00:00:40.05" resultid="5190" heatid="4865" lane="4" entrytime="00:00:41.79" />
                <RESULT eventid="1124" points="212" reactiontime="0" swimtime="00:01:15.15" resultid="5191" heatid="4879" lane="4" entrytime="00:01:17.98" />
                <RESULT eventid="1264" points="213" reactiontime="0" swimtime="00:00:33.75" resultid="5192" heatid="4926" lane="3" entrytime="00:00:36.13" />
                <RESULT eventid="1312" points="153" reactiontime="0" swimtime="00:00:40.58" resultid="5193" heatid="4943" lane="4" entrytime="00:00:41.08" />
                <RESULT eventid="1392" points="167" reactiontime="0" swimtime="00:01:27.76" resultid="5194" heatid="4962" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1420" points="211" reactiontime="0" swimtime="00:02:46.80" resultid="5195" heatid="4969" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                    <SPLIT distance="100" swimtime="00:01:24.39" />
                    <SPLIT distance="150" swimtime="00:02:06.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathan" lastname="Novak Pinho" birthdate="2012-11-14" gender="M" nation="BRA" license="378199" swrid="5603879" athleteid="4410" externalid="378199">
              <RESULTS>
                <RESULT eventid="1096" points="97" reactiontime="0" swimtime="00:00:48.25" resultid="5196" heatid="4865" lane="2" entrytime="00:00:49.68" />
                <RESULT eventid="1124" points="136" reactiontime="0" swimtime="00:01:27.01" resultid="5197" heatid="4878" lane="4" entrytime="00:01:31.09" />
                <RESULT eventid="1264" points="130" reactiontime="0" swimtime="00:00:39.75" resultid="5198" heatid="4925" lane="5" entrytime="00:00:40.86" />
                <RESULT eventid="1392" points="95" reactiontime="0" swimtime="00:01:45.85" resultid="5199" heatid="4962" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1420" points="150" reactiontime="0" swimtime="00:03:06.78" resultid="5200" heatid="4968" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.86" />
                    <SPLIT distance="100" swimtime="00:01:30.13" />
                    <SPLIT distance="150" swimtime="00:02:19.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Antônio Boeing" birthdate="2004-06-04" gender="M" nation="BRA" license="317474" swrid="5184340" athleteid="4240" externalid="317474">
              <RESULTS>
                <RESULT eventid="1075" points="549" reactiontime="0" swimtime="00:02:13.83" resultid="5056" heatid="4856" lane="4" entrytime="00:02:13.88" />
                <RESULT eventid="1135" points="420" reactiontime="0" swimtime="00:00:59.85" resultid="5057" heatid="4885" lane="4" entrytime="00:00:53.87" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Antonio Mendes" birthdate="2008-12-04" gender="M" nation="BRA" license="366962" swrid="5196287" athleteid="4292" externalid="366962">
              <RESULTS>
                <RESULT eventid="1107" points="325" reactiontime="0" swimtime="00:00:32.30" resultid="5097" heatid="4867" lane="3" />
                <RESULT eventid="1183" points="421" reactiontime="0" swimtime="00:00:33.27" resultid="5098" heatid="4900" lane="6" entrytime="00:00:34.54" />
                <RESULT eventid="1243" points="393" reactiontime="0" swimtime="00:02:43.94" resultid="5099" heatid="4912" lane="2" entrytime="00:02:47.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.66" />
                    <SPLIT distance="100" swimtime="00:01:18.19" />
                    <SPLIT distance="150" swimtime="00:02:00.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1377" points="427" reactiontime="0" swimtime="00:01:13.36" resultid="5100" heatid="4960" lane="5" entrytime="00:01:15.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1403" points="281" reactiontime="0" swimtime="00:01:13.70" resultid="5101" heatid="4964" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Camila Cuenca" birthdate="2005-10-06" gender="F" nation="BRA" license="308081" swrid="5357445" athleteid="4243" externalid="308081">
              <RESULTS>
                <RESULT eventid="1127" points="471" reactiontime="0" swimtime="00:01:04.58" resultid="5058" heatid="4881" lane="4" entrytime="00:01:02.48" />
                <RESULT eventid="1267" points="465" reactiontime="0" swimtime="00:00:29.58" resultid="5059" heatid="4928" lane="4" entrytime="00:00:28.49" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Carneiro" birthdate="2010-04-22" gender="F" nation="BRA" license="370670" swrid="5369598" athleteid="4464" externalid="370670">
              <RESULTS>
                <RESULT eventid="1067" points="359" reactiontime="0" swimtime="00:02:51.36" resultid="5241" heatid="4853" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.48" />
                    <SPLIT distance="100" swimtime="00:01:22.86" />
                    <SPLIT distance="150" swimtime="00:02:15.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="427" reactiontime="0" swimtime="00:01:06.72" resultid="5242" heatid="4881" lane="7" entrytime="00:01:08.83" />
                <RESULT eventid="1267" points="402" reactiontime="0" swimtime="00:00:31.06" resultid="5243" heatid="4928" lane="7" entrytime="00:00:31.67" />
                <RESULT eventid="1315" points="348" reactiontime="0" swimtime="00:00:34.66" resultid="5244" heatid="4944" lane="5" entrytime="00:00:34.24" />
                <RESULT eventid="1353" points="430" reactiontime="0" swimtime="00:02:26.11" resultid="5245" heatid="4955" lane="3" entrytime="00:02:31.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                    <SPLIT distance="100" swimtime="00:01:12.57" />
                    <SPLIT distance="150" swimtime="00:01:50.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1445" points="302" reactiontime="0" swimtime="00:01:21.31" resultid="5246" heatid="4974" lane="5" entrytime="00:01:20.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Paiva Boeing" birthdate="2008-01-22" gender="F" nation="BRA" license="318185" swrid="5603884" athleteid="4249" externalid="318185">
              <RESULTS>
                <RESULT eventid="1127" points="425" reactiontime="0" swimtime="00:01:06.82" resultid="5062" heatid="4881" lane="6" entrytime="00:01:07.57" />
                <RESULT eventid="1175" points="400" reactiontime="0" swimtime="00:00:38.75" resultid="5063" heatid="4897" lane="5" entrytime="00:00:42.44" />
                <RESULT eventid="1267" points="440" reactiontime="0" swimtime="00:00:30.13" resultid="5064" heatid="4928" lane="5" entrytime="00:00:30.22" />
                <RESULT eventid="1315" points="386" reactiontime="0" swimtime="00:00:33.46" resultid="5065" heatid="4944" lane="4" entrytime="00:00:33.99" />
                <RESULT eventid="1353" points="416" reactiontime="0" swimtime="00:02:27.68" resultid="5066" heatid="4955" lane="5" entrytime="00:02:29.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                    <SPLIT distance="100" swimtime="00:01:09.91" />
                    <SPLIT distance="150" swimtime="00:01:49.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Naima" lastname="Martins Celestino" birthdate="2004-08-02" gender="F" nation="BRA" license="281995" swrid="5603871" athleteid="4232" externalid="281995">
              <RESULTS>
                <RESULT eventid="1143" points="473" reactiontime="0" swimtime="00:02:33.49" resultid="5050" heatid="4886" lane="4" entrytime="00:02:31.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                    <SPLIT distance="100" swimtime="00:01:14.21" />
                    <SPLIT distance="150" swimtime="00:01:52.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1445" points="585" reactiontime="0" swimtime="00:01:05.25" resultid="5051" heatid="4974" lane="4" entrytime="00:01:04.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniela" lastname="Inoue" birthdate="2008-10-31" gender="F" nation="BRA" license="378348" swrid="5603856" athleteid="4471" externalid="378348">
              <RESULTS>
                <RESULT eventid="1127" points="292" reactiontime="0" swimtime="00:01:15.73" resultid="5247" heatid="4880" lane="2" entrytime="00:01:25.19" />
                <RESULT eventid="1267" points="301" reactiontime="0" swimtime="00:00:34.21" resultid="5248" heatid="4927" lane="6" entrytime="00:00:37.28" />
                <RESULT eventid="1315" points="239" reactiontime="0" swimtime="00:00:39.28" resultid="5249" heatid="4944" lane="7" entrytime="00:00:44.38" />
                <RESULT eventid="1445" points="183" reactiontime="0" swimtime="00:01:36.01" resultid="5250" heatid="4974" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Junio Brambilla" birthdate="2002-04-08" gender="M" nation="BRA" license="392112" swrid="5603859" athleteid="4563" externalid="392112">
              <RESULTS>
                <RESULT eventid="1275" points="270" reactiontime="0" swimtime="00:00:31.16" resultid="5321" heatid="4929" lane="6" />
                <RESULT eventid="1323" points="306" reactiontime="0" swimtime="00:00:32.26" resultid="5322" heatid="4946" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raphael" lastname="Piai Pellegrini" birthdate="2012-03-24" gender="M" nation="BRA" license="377261" swrid="5603894" athleteid="4383" externalid="377261">
              <RESULTS>
                <RESULT eventid="1096" points="143" reactiontime="0" swimtime="00:00:42.49" resultid="5173" heatid="4865" lane="6" entrytime="00:00:47.68" />
                <RESULT eventid="1124" points="179" reactiontime="0" swimtime="00:01:19.45" resultid="5174" heatid="4879" lane="2" entrytime="00:01:24.70" />
                <RESULT eventid="1264" points="198" reactiontime="0" swimtime="00:00:34.54" resultid="5175" heatid="4926" lane="6" entrytime="00:00:36.38" />
                <RESULT eventid="1312" points="119" reactiontime="0" swimtime="00:00:44.12" resultid="5176" heatid="4942" lane="4" entrytime="00:01:02.64" />
                <RESULT eventid="1392" points="126" reactiontime="0" swimtime="00:01:36.34" resultid="5177" heatid="4962" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1420" points="183" reactiontime="0" swimtime="00:02:54.84" resultid="5178" heatid="4969" lane="3" entrytime="00:03:39.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.73" />
                    <SPLIT distance="100" swimtime="00:01:23.81" />
                    <SPLIT distance="150" swimtime="00:02:11.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Carolina Cordeiro" birthdate="2011-04-10" gender="F" nation="BRA" license="392102" swrid="5378340" athleteid="4516" externalid="392102">
              <RESULTS>
                <RESULT eventid="1093" points="36" reactiontime="0" swimtime="00:01:16.13" resultid="5283" heatid="4861" lane="3" />
                <RESULT eventid="1261" points="39" reactiontime="0" swimtime="00:01:07.23" resultid="5284" heatid="4920" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amanda" lastname="Seravalli Zani" birthdate="2014-05-19" gender="F" nation="BRA" license="392096" swrid="5603910" athleteid="4486" externalid="392096">
              <RESULTS>
                <RESULT eventid="1163" points="82" reactiontime="0" swimtime="00:01:05.66" resultid="5259" heatid="4890" lane="7" />
                <RESULT eventid="1255" points="59" reactiontime="0" swimtime="00:00:58.65" resultid="5260" heatid="4915" lane="6" />
                <RESULT eventid="1303" points="48" reactiontime="0" swimtime="00:01:06.91" resultid="5261" heatid="4936" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Quental De Meireles" birthdate="2008-11-20" gender="M" nation="BRA" license="392103" swrid="5603898" athleteid="4519" externalid="392103">
              <RESULTS>
                <RESULT eventid="1135" points="184" reactiontime="0" swimtime="00:01:18.70" resultid="5285" heatid="4882" lane="5" />
                <RESULT eventid="1183" points="168" reactiontime="0" swimtime="00:00:45.15" resultid="5286" heatid="4898" lane="3" />
                <RESULT eventid="1275" points="186" reactiontime="0" swimtime="00:00:35.30" resultid="5287" heatid="4929" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Rampasi" birthdate="2013-10-16" gender="F" nation="BRA" license="382209" swrid="5603866" athleteid="4428" externalid="382209">
              <RESULTS>
                <RESULT eventid="1087" points="68" reactiontime="0" swimtime="00:01:01.77" resultid="5211" heatid="4859" lane="7" entrytime="00:01:05.76" />
                <RESULT eventid="1115" points="98" reactiontime="0" swimtime="00:01:48.95" resultid="5212" heatid="4871" lane="2" entrytime="00:01:55.88" />
                <RESULT eventid="1255" points="100" reactiontime="0" swimtime="00:00:49.31" resultid="5213" heatid="4916" lane="2" entrytime="00:00:52.88" />
                <RESULT eventid="1303" points="46" reactiontime="0" swimtime="00:01:07.76" resultid="5214" heatid="4937" lane="3" entrytime="00:01:11.28" />
                <RESULT eventid="1411" points="111" reactiontime="0" swimtime="00:03:48.93" resultid="5215" heatid="4965" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.65" />
                    <SPLIT distance="100" swimtime="00:01:55.90" />
                    <SPLIT distance="150" swimtime="00:02:55.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Dos Monteiro" birthdate="2014-08-05" gender="M" nation="BRA" license="392095" swrid="5494354" athleteid="4481" externalid="392095">
              <RESULTS>
                <RESULT eventid="1118" points="132" reactiontime="0" swimtime="00:01:28.02" resultid="5255" heatid="4873" lane="2" />
                <RESULT eventid="1166" points="94" reactiontime="0" swimtime="00:00:54.80" resultid="5256" heatid="4892" lane="5" />
                <RESULT eventid="1258" points="125" reactiontime="0" swimtime="00:00:40.23" resultid="5257" heatid="4917" lane="5" />
                <RESULT eventid="1306" points="68" reactiontime="0" swimtime="00:00:53.03" resultid="5258" heatid="4939" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Tomazeli" birthdate="2013-02-05" gender="M" nation="BRA" license="392109" swrid="5614097" athleteid="5308" externalid="392109">
              <RESULTS>
                <RESULT eventid="1090" points="73" reactiontime="0" swimtime="00:00:53.02" resultid="5309" heatid="4860" lane="7" />
                <RESULT eventid="1118" points="56" reactiontime="0" swimtime="00:01:56.79" resultid="5310" heatid="4873" lane="6" />
                <RESULT eventid="1258" points="77" reactiontime="0" swimtime="00:00:47.31" resultid="5311" heatid="4919" lane="7" />
                <RESULT eventid="1306" points="39" reactiontime="0" swimtime="00:01:04.08" resultid="5312" heatid="4938" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Chaim" birthdate="2011-05-29" gender="F" nation="BRA" license="370662" swrid="5409721" athleteid="4351" externalid="370662">
              <RESULTS>
                <RESULT eventid="1061" points="176" reactiontime="0" swimtime="00:03:37.24" resultid="5146" heatid="4850" lane="5" />
                <RESULT eventid="1121" points="220" reactiontime="0" swimtime="00:01:23.15" resultid="5147" heatid="4875" lane="5" entrytime="00:01:26.94" />
                <RESULT eventid="1229" points="227" reactiontime="0" swimtime="00:06:23.30" resultid="5148" heatid="4908" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.16" />
                    <SPLIT distance="100" swimtime="00:01:30.53" />
                    <SPLIT distance="150" swimtime="00:02:20.36" />
                    <SPLIT distance="200" swimtime="00:03:09.26" />
                    <SPLIT distance="250" swimtime="00:03:59.23" />
                    <SPLIT distance="300" swimtime="00:04:48.63" />
                    <SPLIT distance="350" swimtime="00:05:38.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1261" points="229" reactiontime="0" swimtime="00:00:37.43" resultid="5149" heatid="4922" lane="5" entrytime="00:00:38.01" />
                <RESULT eventid="1389" points="161" reactiontime="0" swimtime="00:01:40.80" resultid="5150" heatid="4961" lane="4" entrytime="00:01:47.07" />
                <RESULT eventid="1417" points="194" reactiontime="0" swimtime="00:03:10.50" resultid="5151" heatid="4967" lane="4" entrytime="00:03:02.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.17" />
                    <SPLIT distance="100" swimtime="00:01:31.60" />
                    <SPLIT distance="150" swimtime="00:02:22.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ramon" lastname="Veiga" birthdate="2005-03-31" gender="M" nation="BRA" license="348598" swrid="5603925" athleteid="4264" externalid="348598">
              <RESULTS>
                <RESULT eventid="1135" points="237" reactiontime="0" swimtime="00:01:12.40" resultid="5074" heatid="4882" lane="4" />
                <RESULT eventid="1183" points="442" reactiontime="0" swimtime="00:00:32.73" resultid="5075" heatid="4900" lane="5" entrytime="00:00:32.16" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Marques Picolo" birthdate="2010-07-01" gender="M" nation="BRA" license="366990" swrid="5603869" athleteid="4571" externalid="366990">
              <RESULTS>
                <RESULT eventid="1135" points="211" reactiontime="0" swimtime="00:01:15.31" resultid="5327" heatid="4882" lane="6" />
                <RESULT eventid="1183" reactiontime="0" status="DSQ" swimtime="00:00:00.00" resultid="5328" heatid="4898" lane="4" />
                <RESULT eventid="1275" points="201" reactiontime="0" swimtime="00:00:34.36" resultid="5329" heatid="4929" lane="7" />
                <RESULT eventid="1323" points="119" reactiontime="0" swimtime="00:00:44.12" resultid="5330" heatid="4946" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Hugo Santos" birthdate="2007-03-26" gender="M" nation="BRA" license="384355" swrid="5603855" athleteid="4453" externalid="384355">
              <RESULTS>
                <RESULT eventid="1107" points="185" reactiontime="0" swimtime="00:00:38.94" resultid="5232" heatid="4867" lane="5" />
                <RESULT eventid="1135" points="236" reactiontime="0" swimtime="00:01:12.48" resultid="5233" heatid="4883" lane="4" entrytime="00:01:13.31" />
                <RESULT eventid="1275" points="235" reactiontime="0" swimtime="00:00:32.66" resultid="5234" heatid="4930" lane="4" entrytime="00:00:33.51" />
                <RESULT eventid="1361" points="249" reactiontime="0" swimtime="00:02:37.79" resultid="5235" heatid="4956" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="100" swimtime="00:01:13.04" />
                    <SPLIT distance="150" swimtime="00:01:55.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Gabriel Oliveira" birthdate="2006-05-31" gender="M" nation="BRA" license="345589" swrid="5603838" athleteid="4312" externalid="345589">
              <RESULTS>
                <RESULT eventid="1135" points="395" reactiontime="0" swimtime="00:01:01.09" resultid="5114" heatid="4884" lane="3" entrytime="00:01:04.52" />
                <RESULT eventid="1275" points="381" reactiontime="0" swimtime="00:00:27.79" resultid="5115" heatid="4931" lane="4" entrytime="00:00:29.29" />
                <RESULT eventid="1323" points="305" reactiontime="0" swimtime="00:00:32.29" resultid="5116" heatid="4946" lane="3" entrytime="00:00:55.68" />
                <RESULT eventid="1361" points="343" reactiontime="0" swimtime="00:02:21.92" resultid="5117" heatid="4956" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                    <SPLIT distance="100" swimtime="00:01:08.12" />
                    <SPLIT distance="150" swimtime="00:01:45.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tiago" lastname="Ficher Delmont Pais" birthdate="2010-07-15" gender="M" nation="BRA" license="338533" swrid="5588701" athleteid="4305" externalid="338533">
              <RESULTS>
                <RESULT eventid="1075" points="355" reactiontime="0" swimtime="00:02:34.77" resultid="5108" heatid="4856" lane="2" entrytime="00:02:37.51" />
                <RESULT eventid="1151" points="317" reactiontime="0" swimtime="00:02:38.62" resultid="5109" heatid="4887" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:18.24" />
                    <SPLIT distance="100" swimtime="00:02:00.36" />
                    <SPLIT distance="150" swimtime="00:02:40.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1291" points="327" reactiontime="0" swimtime="00:02:33.23" resultid="5110" heatid="4934" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.84" />
                    <SPLIT distance="100" swimtime="00:01:14.04" />
                    <SPLIT distance="150" swimtime="00:01:53.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1339" reactiontime="0" status="DSQ" swimtime="00:00:00.00" resultid="5111" heatid="4949" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                    <SPLIT distance="100" swimtime="00:01:11.79" />
                    <SPLIT distance="150" swimtime="00:01:55.91" />
                    <SPLIT distance="200" swimtime="00:02:38.76" />
                    <SPLIT distance="250" swimtime="00:03:26.00" />
                    <SPLIT distance="300" swimtime="00:04:14.50" />
                    <SPLIT distance="350" swimtime="00:04:53.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" points="391" reactiontime="0" swimtime="00:02:15.79" resultid="5112" heatid="4957" lane="2" entrytime="00:02:17.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                    <SPLIT distance="100" swimtime="00:01:05.73" />
                    <SPLIT distance="150" swimtime="00:01:40.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" points="375" reactiontime="0" swimtime="00:01:06.25" resultid="5113" heatid="4975" lane="4" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Corsine Ferreira" birthdate="2010-03-10" gender="F" nation="BRA" license="353591" swrid="5588608" athleteid="4458" externalid="353591">
              <RESULTS>
                <RESULT eventid="1067" points="313" reactiontime="0" swimtime="00:02:59.34" resultid="5236" heatid="4853" lane="4" entrytime="00:02:59.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.93" />
                    <SPLIT distance="100" swimtime="00:01:23.44" />
                    <SPLIT distance="150" swimtime="00:02:17.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="320" reactiontime="0" swimtime="00:11:40.29" resultid="5237" heatid="4901" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:11:42.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1283" points="375" reactiontime="0" swimtime="00:02:44.82" resultid="5238" heatid="4933" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.61" />
                    <SPLIT distance="100" swimtime="00:01:20.99" />
                    <SPLIT distance="150" swimtime="00:02:03.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1353" points="326" reactiontime="0" swimtime="00:02:40.27" resultid="5239" heatid="4955" lane="6" entrytime="00:02:37.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                    <SPLIT distance="100" swimtime="00:01:16.67" />
                    <SPLIT distance="150" swimtime="00:01:58.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1395" points="350" reactiontime="0" swimtime="00:01:17.88" resultid="5240" heatid="4963" lane="5" entrytime="00:01:19.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Henrique Goes" birthdate="2008-10-26" gender="M" nation="BRA" license="392105" swrid="5603853" athleteid="4527" externalid="392105">
              <RESULTS>
                <RESULT eventid="1075" points="159" reactiontime="0" swimtime="00:03:22.11" resultid="5291" heatid="4855" lane="6" />
                <RESULT eventid="1183" points="136" reactiontime="0" swimtime="00:00:48.49" resultid="5292" heatid="4899" lane="2" />
                <RESULT eventid="1275" points="160" reactiontime="0" swimtime="00:00:37.07" resultid="5293" heatid="4929" lane="3" />
                <RESULT eventid="1323" points="98" reactiontime="0" swimtime="00:00:47.16" resultid="5294" heatid="4945" lane="4" />
                <RESULT eventid="1377" points="149" reactiontime="0" swimtime="00:01:44.17" resultid="5295" heatid="4959" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Furuchi Martins" birthdate="2011-10-05" gender="F" nation="BRA" license="367001" swrid="5602616" athleteid="4566" externalid="367001">
              <RESULTS>
                <RESULT eventid="1121" points="122" reactiontime="0" swimtime="00:01:41.05" resultid="5323" heatid="4874" lane="5" />
                <RESULT eventid="1169" points="136" reactiontime="0" swimtime="00:00:55.43" resultid="5324" heatid="4893" lane="3" />
                <RESULT eventid="1261" points="157" reactiontime="0" swimtime="00:00:42.44" resultid="5325" heatid="4920" lane="6" />
                <RESULT eventid="1347" points="153" reactiontime="0" swimtime="00:01:56.39" resultid="5326" heatid="4950" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernando" lastname="Santin Dolis" birthdate="2008-12-18" gender="M" nation="BRA" license="355590" swrid="5603907" athleteid="4255" externalid="355590">
              <RESULTS>
                <RESULT eventid="1075" points="204" reactiontime="0" swimtime="00:03:06.01" resultid="5067" heatid="4855" lane="5" entrytime="00:03:02.39" />
                <RESULT eventid="1291" points="192" reactiontime="0" swimtime="00:03:02.80" resultid="5068" heatid="4934" lane="4" entrytime="00:02:48.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.25" />
                    <SPLIT distance="100" swimtime="00:01:27.76" />
                    <SPLIT distance="150" swimtime="00:02:15.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1403" points="206" reactiontime="0" swimtime="00:01:21.73" resultid="5069" heatid="4964" lane="5" entrytime="00:01:20.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Bessa" birthdate="2003-06-19" gender="M" nation="BRA" license="317841" swrid="5312237" athleteid="4206" externalid="317841">
              <RESULTS>
                <RESULT eventid="1135" points="491" reactiontime="0" swimtime="00:00:56.83" resultid="5029" heatid="4885" lane="6" entrytime="00:00:57.78" />
                <RESULT eventid="1243" points="588" reactiontime="0" swimtime="00:02:23.41" resultid="5030" heatid="4912" lane="4" entrytime="00:02:22.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                    <SPLIT distance="100" swimtime="00:01:09.48" />
                    <SPLIT distance="150" swimtime="00:01:45.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Sol Reolon Gomes" birthdate="2011-02-28" gender="F" nation="BRA" license="392100" swrid="5603914" athleteid="4506" externalid="392100">
              <RESULTS>
                <RESULT eventid="1093" points="141" reactiontime="0" swimtime="00:00:48.51" resultid="5275" heatid="4861" lane="7" />
                <RESULT eventid="1121" points="165" reactiontime="0" swimtime="00:01:31.44" resultid="5276" heatid="4874" lane="3" />
                <RESULT eventid="1261" points="198" reactiontime="0" swimtime="00:00:39.34" resultid="5277" heatid="4921" lane="7" />
                <RESULT eventid="1309" points="118" reactiontime="0" swimtime="00:00:49.60" resultid="5278" heatid="4940" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lara" lastname="Constantino" birthdate="2012-06-02" gender="F" nation="BRA" license="382208" swrid="5420069" athleteid="4422" externalid="382208">
              <RESULTS>
                <RESULT eventid="1121" points="164" reactiontime="0" swimtime="00:01:31.68" resultid="5206" heatid="4875" lane="3" entrytime="00:01:34.58" />
                <RESULT eventid="1169" points="203" reactiontime="0" swimtime="00:00:48.55" resultid="5207" heatid="4894" lane="5" entrytime="00:00:50.37" />
                <RESULT eventid="1261" points="181" reactiontime="0" swimtime="00:00:40.50" resultid="5208" heatid="4922" lane="3" entrytime="00:00:40.88" />
                <RESULT eventid="1347" points="181" reactiontime="0" swimtime="00:01:50.14" resultid="5209" heatid="4951" lane="6" />
                <RESULT eventid="1417" points="143" reactiontime="0" swimtime="00:03:30.80" resultid="5210" heatid="4967" lane="3" entrytime="00:03:33.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.87" />
                    <SPLIT distance="100" swimtime="00:01:45.73" />
                    <SPLIT distance="150" swimtime="00:02:41.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Otavio Costa" birthdate="2009-01-28" gender="M" nation="BRA" license="370666" swrid="5603881" athleteid="4364" externalid="370666">
              <RESULTS>
                <RESULT eventid="1075" points="176" reactiontime="0" swimtime="00:03:15.45" resultid="5157" heatid="4855" lane="3" />
                <RESULT eventid="1135" points="189" reactiontime="0" swimtime="00:01:18.11" resultid="5158" heatid="4883" lane="7" />
                <RESULT eventid="1275" points="198" reactiontime="0" swimtime="00:00:34.54" resultid="5159" heatid="4929" lane="5" entrytime="00:00:42.12" />
                <RESULT eventid="1323" points="153" reactiontime="0" swimtime="00:00:40.63" resultid="5160" heatid="4946" lane="5" entrytime="00:00:41.38" />
                <RESULT eventid="1377" points="186" reactiontime="0" swimtime="00:01:36.80" resultid="5161" heatid="4960" lane="2" entrytime="00:01:38.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1453" reactiontime="0" status="DSQ" swimtime="00:00:00.00" resultid="5162" heatid="4975" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Otavio Luz" birthdate="2013-07-27" gender="M" nation="BRA" license="392111" swrid="5603882" athleteid="4558" externalid="392111">
              <RESULTS>
                <RESULT eventid="1118" points="93" reactiontime="0" swimtime="00:01:38.89" resultid="5317" heatid="4872" lane="6" />
                <RESULT eventid="1166" points="40" reactiontime="0" swimtime="00:01:12.42" resultid="5318" heatid="4891" lane="4" />
                <RESULT eventid="1258" points="103" reactiontime="0" swimtime="00:00:43.00" resultid="5319" heatid="4917" lane="4" />
                <RESULT eventid="1306" points="38" reactiontime="0" swimtime="00:01:04.19" resultid="5320" heatid="4939" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Assuncao Silva" birthdate="2012-11-11" gender="M" nation="BRA" license="392110" swrid="5200167" athleteid="4553" externalid="392110">
              <RESULTS>
                <RESULT eventid="1124" points="130" reactiontime="0" swimtime="00:01:28.45" resultid="5313" heatid="4877" lane="7" />
                <RESULT eventid="1172" points="124" reactiontime="0" swimtime="00:00:49.93" resultid="5314" heatid="4895" lane="6" />
                <RESULT eventid="1264" points="142" reactiontime="0" swimtime="00:00:38.57" resultid="5315" heatid="4923" lane="5" />
                <RESULT eventid="1350" points="118" reactiontime="0" swimtime="00:01:52.69" resultid="5316" heatid="4953" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robsson" lastname="Tows Oliveira" birthdate="2014-03-05" gender="M" nation="BRA" license="392107" swrid="5603922" athleteid="4538" externalid="392107">
              <RESULTS>
                <RESULT eventid="1118" points="94" reactiontime="0" swimtime="00:01:38.35" resultid="5300" heatid="4873" lane="7" />
                <RESULT eventid="1166" points="98" reactiontime="0" swimtime="00:00:53.94" resultid="5301" heatid="4891" lane="3" />
                <RESULT eventid="1210" points="84" reactiontime="0" swimtime="00:01:52.42" resultid="5302" heatid="4905" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="95" reactiontime="0" swimtime="00:00:44.16" resultid="5303" heatid="4918" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Sanches Ghelere" birthdate="2008-08-06" gender="F" nation="BRA" license="372024" swrid="5603905" athleteid="4286" externalid="372024">
              <RESULTS>
                <RESULT eventid="1127" points="458" reactiontime="0" swimtime="00:01:05.15" resultid="5092" heatid="4881" lane="2" entrytime="00:01:08.56" />
                <RESULT eventid="1191" points="381" reactiontime="0" swimtime="00:11:00.66" resultid="5093" heatid="4901" lane="6" />
                <RESULT eventid="1267" points="457" reactiontime="0" swimtime="00:00:29.76" resultid="5094" heatid="4928" lane="6" entrytime="00:00:30.49" />
                <RESULT eventid="1315" points="418" reactiontime="0" swimtime="00:00:32.60" resultid="5095" heatid="4944" lane="3" entrytime="00:00:34.54" />
                <RESULT eventid="1445" points="407" reactiontime="0" swimtime="00:01:13.62" resultid="5096" heatid="4974" lane="3" entrytime="00:01:22.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Garcia Cavalcante" birthdate="2011-11-21" gender="M" nation="BRA" license="378200" swrid="5603840" athleteid="4416" externalid="378200">
              <RESULTS>
                <RESULT eventid="1124" points="176" reactiontime="0" swimtime="00:01:19.88" resultid="5201" heatid="4879" lane="7" entrytime="00:01:26.07" />
                <RESULT eventid="1172" points="192" reactiontime="0" swimtime="00:00:43.18" resultid="5202" heatid="4896" lane="5" entrytime="00:00:47.20" />
                <RESULT eventid="1264" points="179" reactiontime="0" swimtime="00:00:35.76" resultid="5203" heatid="4926" lane="2" entrytime="00:00:38.46" />
                <RESULT eventid="1350" points="174" reactiontime="0" swimtime="00:01:38.93" resultid="5204" heatid="4953" lane="5" entrytime="00:01:45.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1420" points="174" reactiontime="0" swimtime="00:02:57.75" resultid="5205" heatid="4969" lane="5" entrytime="00:03:13.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.99" />
                    <SPLIT distance="100" swimtime="00:01:26.95" />
                    <SPLIT distance="150" swimtime="00:02:15.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Borges Carneiro" birthdate="1998-05-07" gender="F" nation="BRA" license="266382" swrid="5339063" athleteid="4235" externalid="266382">
              <RESULTS>
                <RESULT eventid="1127" points="483" reactiontime="0" swimtime="00:01:04.01" resultid="5052" heatid="4881" lane="3" entrytime="00:01:03.96" />
                <RESULT eventid="1175" points="578" reactiontime="0" swimtime="00:00:34.28" resultid="5053" heatid="4897" lane="4" entrytime="00:00:36.00" />
                <RESULT eventid="1331" points="416" reactiontime="0" swimtime="00:05:46.68" resultid="5054" heatid="4948" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                    <SPLIT distance="100" swimtime="00:01:19.57" />
                    <SPLIT distance="150" swimtime="00:02:07.89" />
                    <SPLIT distance="200" swimtime="00:02:54.03" />
                    <SPLIT distance="250" swimtime="00:03:38.44" />
                    <SPLIT distance="300" swimtime="00:04:24.97" />
                    <SPLIT distance="350" swimtime="00:05:06.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1369" points="532" reactiontime="0" swimtime="00:01:16.94" resultid="5055" heatid="4958" lane="4" entrytime="00:01:17.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Osmar" lastname="Campos" birthdate="2012-06-04" gender="M" nation="BRA" license="377264" swrid="5362294" athleteid="4396" externalid="377264">
              <RESULTS>
                <RESULT eventid="1096" points="107" reactiontime="0" swimtime="00:00:46.73" resultid="5184" heatid="4864" lane="4" entrytime="00:00:55.39" />
                <RESULT eventid="1124" points="134" reactiontime="0" swimtime="00:01:27.58" resultid="5185" heatid="4878" lane="3" entrytime="00:01:41.38" />
                <RESULT eventid="1264" points="139" reactiontime="0" swimtime="00:00:38.84" resultid="5186" heatid="4925" lane="2" entrytime="00:00:45.11" />
                <RESULT eventid="1312" points="67" reactiontime="0" swimtime="00:00:53.39" resultid="5187" heatid="4943" lane="6" entrytime="00:00:58.88" />
                <RESULT eventid="1420" points="147" reactiontime="0" swimtime="00:03:08.15" resultid="5188" heatid="4968" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.29" />
                    <SPLIT distance="100" swimtime="00:01:31.01" />
                    <SPLIT distance="150" swimtime="00:02:20.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1442" points="57" reactiontime="0" swimtime="00:02:03.74" resultid="5189" heatid="4973" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Batista Sanchez" birthdate="2009-05-22" gender="M" nation="BRA" license="370668" swrid="5255779" athleteid="4221" externalid="370668">
              <RESULTS>
                <RESULT eventid="1183" points="309" reactiontime="0" swimtime="00:00:36.89" resultid="5041" heatid="4900" lane="2" entrytime="00:00:40.13" />
                <RESULT eventid="1243" points="289" reactiontime="0" swimtime="00:03:01.61" resultid="5042" heatid="4911" lane="5" entrytime="00:03:05.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                    <SPLIT distance="100" swimtime="00:01:25.51" />
                    <SPLIT distance="150" swimtime="00:02:13.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1323" points="229" reactiontime="0" swimtime="00:00:35.53" resultid="5043" heatid="4946" lane="6" />
                <RESULT eventid="1377" points="307" reactiontime="0" swimtime="00:01:21.94" resultid="5044" heatid="4960" lane="6" entrytime="00:01:26.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1431" points="210" reactiontime="0" swimtime="00:01:22.90" resultid="5045" heatid="4971" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felype" lastname="Gongora Zago" birthdate="2011-09-14" gender="M" nation="BRA" license="392099" swrid="5603848" athleteid="4501" externalid="392099">
              <RESULTS>
                <RESULT eventid="1096" points="79" reactiontime="0" swimtime="00:00:51.70" resultid="5271" heatid="4864" lane="5" />
                <RESULT eventid="1124" points="75" reactiontime="0" swimtime="00:01:46.23" resultid="5272" heatid="4876" lane="5" />
                <RESULT eventid="1264" points="72" reactiontime="0" swimtime="00:00:48.31" resultid="5273" heatid="4923" lane="6" />
                <RESULT eventid="1392" reactiontime="0" status="DSQ" swimtime="00:00:00.00" resultid="5274" heatid="4962" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otavio" lastname="Sossai Altoé" birthdate="2006-09-04" gender="M" nation="BRA" license="296488" swrid="5603915" athleteid="4202" externalid="296488">
              <RESULTS>
                <RESULT eventid="1135" points="585" reactiontime="0" swimtime="00:00:53.60" resultid="5026" heatid="4885" lane="5" entrytime="00:00:54.70" />
                <RESULT eventid="1275" points="512" reactiontime="0" swimtime="00:00:25.19" resultid="5027" heatid="4932" lane="4" entrytime="00:00:25.16" />
                <RESULT eventid="1361" points="594" reactiontime="0" swimtime="00:01:58.18" resultid="5028" heatid="4957" lane="4" entrytime="00:01:59.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.51" />
                    <SPLIT distance="100" swimtime="00:00:56.01" />
                    <SPLIT distance="150" swimtime="00:01:26.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Diogo" lastname="Sanchez" birthdate="2012-11-29" gender="M" nation="BRA" license="370658" swrid="5603906" athleteid="4340" externalid="370658">
              <RESULTS>
                <RESULT eventid="1124" points="65" reactiontime="0" swimtime="00:01:51.00" resultid="5137" heatid="4877" lane="4" entrytime="00:02:00.64" />
                <RESULT eventid="1172" points="73" reactiontime="0" swimtime="00:00:59.62" resultid="5138" heatid="4896" lane="7" entrytime="00:01:01.56" />
                <RESULT eventid="1264" points="66" reactiontime="0" swimtime="00:00:49.69" resultid="5139" heatid="4924" lane="4" entrytime="00:00:54.74" />
                <RESULT eventid="1350" points="66" reactiontime="0" swimtime="00:02:16.18" resultid="5140" heatid="4952" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietro" lastname="Nabas De Assis" birthdate="2011-07-09" gender="M" nation="BRA" license="366968" swrid="5603878" athleteid="4327" externalid="366968">
              <RESULTS>
                <RESULT eventid="1064" points="166" reactiontime="0" swimtime="00:03:19.43" resultid="5126" heatid="4852" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.93" />
                    <SPLIT distance="100" swimtime="00:01:37.24" />
                    <SPLIT distance="150" swimtime="00:02:33.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="173" reactiontime="0" swimtime="00:00:44.71" resultid="5127" heatid="4896" lane="4" entrytime="00:00:44.96" />
                <RESULT eventid="1264" points="175" reactiontime="0" swimtime="00:00:36.00" resultid="5128" heatid="4926" lane="5" entrytime="00:00:35.86" />
                <RESULT eventid="1350" points="144" reactiontime="0" swimtime="00:01:45.37" resultid="5129" heatid="4953" lane="4" entrytime="00:01:41.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1420" points="196" reactiontime="0" swimtime="00:02:50.88" resultid="5130" heatid="4969" lane="4" entrytime="00:02:51.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                    <SPLIT distance="100" swimtime="00:01:20.82" />
                    <SPLIT distance="150" swimtime="00:02:06.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caetano" lastname="Alves Santos" birthdate="2013-09-03" gender="M" nation="BRA" license="392101" swrid="5179765" athleteid="4511" externalid="392101">
              <RESULTS>
                <RESULT eventid="1118" points="65" reactiontime="0" swimtime="00:01:51.03" resultid="5279" heatid="4873" lane="3" />
                <RESULT eventid="1166" points="41" reactiontime="0" swimtime="00:01:12.32" resultid="5280" heatid="4892" lane="3" />
                <RESULT eventid="1258" points="70" reactiontime="0" swimtime="00:00:48.78" resultid="5281" heatid="4918" lane="2" />
                <RESULT eventid="1306" points="26" reactiontime="0" swimtime="00:01:13.28" resultid="5282" heatid="4938" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Garcia Cavalcante" birthdate="2008-08-11" gender="M" nation="BRA" license="369676" swrid="5603841" athleteid="4227" externalid="369676">
              <RESULTS>
                <RESULT eventid="1075" points="313" reactiontime="0" swimtime="00:02:41.33" resultid="5046" heatid="4855" lane="4" entrytime="00:02:49.87" />
                <RESULT eventid="1243" points="376" reactiontime="0" swimtime="00:02:46.46" resultid="5047" heatid="4912" lane="6" entrytime="00:02:47.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                    <SPLIT distance="100" swimtime="00:01:19.20" />
                    <SPLIT distance="150" swimtime="00:02:02.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1339" points="291" reactiontime="0" swimtime="00:05:54.11" resultid="5048" heatid="4949" lane="3" entrytime="00:05:50.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.07" />
                    <SPLIT distance="100" swimtime="00:01:27.26" />
                    <SPLIT distance="150" swimtime="00:02:17.98" />
                    <SPLIT distance="200" swimtime="00:03:07.13" />
                    <SPLIT distance="250" swimtime="00:03:49.97" />
                    <SPLIT distance="300" swimtime="00:04:33.87" />
                    <SPLIT distance="350" swimtime="00:05:14.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1377" points="371" reactiontime="0" swimtime="00:01:16.91" resultid="5049" heatid="4960" lane="3" entrytime="00:01:18.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Souza" birthdate="2013-09-11" gender="M" nation="BRA" license="382211" swrid="5603916" athleteid="4441" externalid="382211">
              <RESULTS>
                <RESULT eventid="1118" points="127" reactiontime="0" swimtime="00:01:29.19" resultid="5222" heatid="4873" lane="5" entrytime="00:01:51.76" />
                <RESULT eventid="1166" points="72" reactiontime="0" swimtime="00:00:59.78" resultid="5223" heatid="4892" lane="4" entrytime="00:01:07.43" />
                <RESULT eventid="1258" points="123" reactiontime="0" swimtime="00:00:40.43" resultid="5224" heatid="4919" lane="5" entrytime="00:00:48.10" />
                <RESULT eventid="1306" points="62" reactiontime="0" swimtime="00:00:54.95" resultid="5225" heatid="4939" lane="5" />
                <RESULT eventid="1414" points="144" reactiontime="0" swimtime="00:03:09.23" resultid="5226" heatid="4966" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.06" />
                    <SPLIT distance="100" swimtime="00:01:31.76" />
                    <SPLIT distance="150" swimtime="00:02:21.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Ghelere" birthdate="2011-04-03" gender="F" nation="BRA" license="368146" swrid="5603843" athleteid="4333" externalid="368146">
              <RESULTS>
                <RESULT eventid="1061" points="210" reactiontime="0" swimtime="00:03:24.93" resultid="5131" heatid="4851" lane="4" entrytime="00:03:40.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:03:24.93" />
                    <SPLIT distance="100" swimtime="00:03:37.39" />
                    <SPLIT distance="150" swimtime="00:03:37.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="243" reactiontime="0" swimtime="00:01:20.49" resultid="5132" heatid="4875" lane="4" entrytime="00:01:24.31" />
                <RESULT eventid="1261" points="253" reactiontime="0" swimtime="00:00:36.21" resultid="5133" heatid="4922" lane="4" entrytime="00:00:37.60" />
                <RESULT eventid="1309" points="186" reactiontime="0" swimtime="00:00:42.65" resultid="5134" heatid="4941" lane="4" entrytime="00:00:43.49" />
                <RESULT eventid="1417" points="246" reactiontime="0" swimtime="00:02:55.93" resultid="5135" heatid="4967" lane="5" entrytime="00:03:29.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.79" />
                    <SPLIT distance="100" swimtime="00:01:26.45" />
                    <SPLIT distance="150" swimtime="00:02:11.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1439" points="139" reactiontime="0" swimtime="00:01:45.33" resultid="5136" heatid="4972" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Pacheco" birthdate="2012-10-03" gender="M" nation="BRA" license="370663" swrid="5603883" athleteid="4358" externalid="370663">
              <RESULTS>
                <RESULT eventid="1124" points="178" reactiontime="0" swimtime="00:01:19.68" resultid="5152" heatid="4879" lane="3" entrytime="00:01:23.57" />
                <RESULT eventid="1172" points="125" reactiontime="0" swimtime="00:00:49.83" resultid="5153" heatid="4896" lane="3" entrytime="00:00:52.06" />
                <RESULT eventid="1264" points="179" reactiontime="0" swimtime="00:00:35.73" resultid="5154" heatid="4926" lane="7" entrytime="00:00:38.96" />
                <RESULT eventid="1312" points="122" reactiontime="0" swimtime="00:00:43.84" resultid="5155" heatid="4943" lane="5" entrytime="00:00:45.65" />
                <RESULT eventid="1420" points="180" reactiontime="0" swimtime="00:02:55.94" resultid="5156" heatid="4969" lane="6" entrytime="00:03:44.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.51" />
                    <SPLIT distance="100" swimtime="00:01:25.13" />
                    <SPLIT distance="150" swimtime="00:02:13.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Passafaro" birthdate="2009-02-01" gender="F" nation="BRA" license="370673" swrid="5603885" athleteid="4280" externalid="370673">
              <RESULTS>
                <RESULT eventid="1127" points="354" reactiontime="0" swimtime="00:01:10.98" resultid="5087" heatid="4880" lane="4" entrytime="00:01:10.48" />
                <RESULT eventid="1267" points="382" reactiontime="0" swimtime="00:00:31.60" resultid="5088" heatid="4928" lane="2" entrytime="00:00:31.38" />
                <RESULT eventid="1315" points="264" reactiontime="0" swimtime="00:00:37.96" resultid="5089" heatid="4944" lane="6" entrytime="00:00:36.59" />
                <RESULT eventid="1353" points="348" reactiontime="0" swimtime="00:02:36.71" resultid="5090" heatid="4954" lane="4" entrytime="00:02:44.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.49" />
                    <SPLIT distance="100" swimtime="00:01:15.46" />
                    <SPLIT distance="150" swimtime="00:01:56.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1395" points="203" reactiontime="0" swimtime="00:01:33.33" resultid="5091" heatid="4963" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Casavechia Carraro" birthdate="2009-07-28" gender="M" nation="BRA" license="368150" swrid="5384752" athleteid="4267" externalid="368150">
              <RESULTS>
                <RESULT eventid="1135" points="491" reactiontime="0" swimtime="00:00:56.83" resultid="5076" heatid="4885" lane="7" entrytime="00:00:57.96" />
                <RESULT eventid="1199" points="401" reactiontime="0" swimtime="00:19:07.65" resultid="5077" heatid="4902" lane="4" entrytime="00:19:16.12" />
                <RESULT eventid="1221" points="477" reactiontime="0" swimtime="00:04:31.51" resultid="5078" heatid="4907" lane="4" entrytime="00:04:40.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                    <SPLIT distance="100" swimtime="00:01:04.15" />
                    <SPLIT distance="150" swimtime="00:01:38.12" />
                    <SPLIT distance="200" swimtime="00:02:13.05" />
                    <SPLIT distance="250" swimtime="00:02:48.25" />
                    <SPLIT distance="300" swimtime="00:03:23.83" />
                    <SPLIT distance="350" swimtime="00:03:58.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1339" points="313" reactiontime="0" swimtime="00:05:45.79" resultid="5079" heatid="4949" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                    <SPLIT distance="100" swimtime="00:01:12.90" />
                    <SPLIT distance="150" swimtime="00:02:00.61" />
                    <SPLIT distance="200" swimtime="00:02:46.60" />
                    <SPLIT distance="250" swimtime="00:03:37.62" />
                    <SPLIT distance="300" swimtime="00:04:29.19" />
                    <SPLIT distance="350" swimtime="00:05:08.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1361" points="478" reactiontime="0" swimtime="00:02:07.08" resultid="5080" heatid="4957" lane="3" entrytime="00:02:09.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.75" />
                    <SPLIT distance="100" swimtime="00:01:00.21" />
                    <SPLIT distance="150" swimtime="00:01:33.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1469" points="414" reactiontime="0" swimtime="00:09:54.64" resultid="5081" heatid="4977" lane="4" entrytime="00:09:58.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:09:54.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="1035" nation="BRA" clubid="4778" swrid="93778" name="Fundação de Esportes de Campo Mourão" shortname="Fecam">
          <ATHLETES>
            <ATHLETE firstname="Rafael" lastname="Franco Santos" birthdate="2002-01-03" gender="M" nation="BRA" license="290441" swrid="5546064" athleteid="4782" externalid="290441">
              <RESULTS>
                <RESULT eventid="1075" points="338" reactiontime="0" swimtime="00:02:37.23" resultid="5491" heatid="4856" lane="7" entrytime="00:02:39.80" />
                <RESULT eventid="1275" points="480" reactiontime="0" swimtime="00:00:25.74" resultid="5492" heatid="4932" lane="3" entrytime="00:00:25.86" />
                <RESULT eventid="1323" points="459" reactiontime="0" swimtime="00:00:28.18" resultid="5493" heatid="4947" lane="4" entrytime="00:00:28.12" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Osvaldo" lastname="Valarini" birthdate="1988-06-06" gender="M" nation="BRA" license="189703" swrid="5603923" athleteid="4842" externalid="189703">
              <RESULTS>
                <RESULT eventid="1183" points="279" reactiontime="0" swimtime="00:00:38.17" resultid="5534" heatid="4898" lane="5" />
                <RESULT eventid="1243" reactiontime="0" status="DNS" swimtime="00:00:00.00" resultid="5535" />
                <RESULT eventid="1377" points="258" reactiontime="0" swimtime="00:01:26.82" resultid="5536" heatid="4959" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Corassari Boas" birthdate="2012-02-09" gender="F" nation="BRA" license="392158" swrid="5443189" athleteid="4830" externalid="392158">
              <RESULTS>
                <RESULT eventid="1093" reactiontime="0" status="DSQ" swimtime="00:00:00.00" resultid="5526" heatid="4861" lane="6" />
                <RESULT eventid="1261" points="116" reactiontime="0" swimtime="00:00:46.94" resultid="5527" heatid="4920" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaue" lastname="Guilherme Chagas" birthdate="2005-06-29" gender="M" nation="BRA" license="378464" swrid="5603851" athleteid="4805" externalid="378464">
              <RESULTS>
                <RESULT eventid="1135" points="258" reactiontime="0" swimtime="00:01:10.36" resultid="5516" heatid="4883" lane="6" entrytime="00:01:16.81" />
                <RESULT eventid="1275" points="241" reactiontime="0" swimtime="00:00:32.37" resultid="5517" heatid="4930" lane="5" entrytime="00:00:34.37" />
                <RESULT eventid="1323" points="241" reactiontime="0" swimtime="00:00:34.94" resultid="5518" heatid="4947" lane="7" entrytime="00:00:37.20" />
                <RESULT eventid="1361" points="252" reactiontime="0" swimtime="00:02:37.20" resultid="5519" heatid="4956" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                    <SPLIT distance="100" swimtime="00:01:13.23" />
                    <SPLIT distance="150" swimtime="00:01:55.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Keirrison" lastname="Leite Silva" birthdate="2011-08-02" gender="M" nation="BRA" license="392161" swrid="5603864" athleteid="4839" externalid="392161">
              <RESULTS>
                <RESULT eventid="1096" points="62" reactiontime="0" swimtime="00:00:56.10" resultid="5532" heatid="4864" lane="6" />
                <RESULT eventid="1264" points="69" reactiontime="0" swimtime="00:00:49.09" resultid="5533" heatid="4924" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Pedroso Silverio" birthdate="1994-11-21" gender="M" nation="BRA" license="115715" swrid="5603892" athleteid="4779" externalid="115715">
              <RESULTS>
                <RESULT eventid="1199" points="328" reactiontime="0" swimtime="00:20:27.76" resultid="5489" heatid="4902" lane="5" entrytime="00:20:48.09" />
                <RESULT eventid="1221" reactiontime="0" status="DNS" swimtime="00:00:00.00" resultid="5490" entrytime="00:04:55.46" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Ferreira Batista" birthdate="2012-03-29" gender="F" nation="BRA" license="385779" swrid="5532525" athleteid="4813" externalid="385779">
              <RESULTS>
                <RESULT eventid="1093" points="111" reactiontime="0" swimtime="00:00:52.56" resultid="5522" heatid="4862" lane="2" />
                <RESULT eventid="1261" points="103" reactiontime="0" swimtime="00:00:48.81" resultid="5523" heatid="4921" lane="3" entrytime="00:00:55.14" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Batinga Ponchielli" birthdate="2007-01-18" gender="M" nation="BRA" license="378461" swrid="5251143" athleteid="4798" externalid="378461">
              <RESULTS>
                <RESULT eventid="1107" points="234" reactiontime="0" swimtime="00:00:36.01" resultid="5511" heatid="4868" lane="6" entrytime="00:00:39.71" />
                <RESULT eventid="1275" points="261" reactiontime="0" swimtime="00:00:31.54" resultid="5512" heatid="4930" lane="3" entrytime="00:00:34.42" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Franca Rebollo" birthdate="2012-09-26" gender="M" nation="BRA" license="385780" swrid="5538081" athleteid="4816" externalid="385780">
              <RESULTS>
                <RESULT eventid="1096" points="36" reactiontime="0" swimtime="00:01:06.75" resultid="5524" heatid="4864" lane="3" />
                <RESULT eventid="1264" points="46" reactiontime="0" swimtime="00:00:56.24" resultid="5525" heatid="4924" lane="6" entrytime="00:01:04.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Stipp Silva" birthdate="2009-12-02" gender="M" nation="BRA" license="378462" swrid="5603918" athleteid="4801" externalid="378462">
              <RESULTS>
                <RESULT eventid="1135" points="257" reactiontime="0" swimtime="00:01:10.45" resultid="5513" heatid="4883" lane="2" entrytime="00:01:22.11" />
                <RESULT eventid="1183" points="188" reactiontime="0" swimtime="00:00:43.55" resultid="5514" heatid="4899" lane="3" entrytime="00:00:48.47" />
                <RESULT eventid="1275" points="263" reactiontime="0" swimtime="00:00:31.45" resultid="5515" heatid="4930" lane="7" entrytime="00:00:36.15" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Gomes De Souza" birthdate="2006-01-30" gender="F" nation="BRA" license="308464" swrid="5603844" athleteid="4819" externalid="308464">
              <RESULTS>
                <RESULT eventid="1099" points="216" reactiontime="0" swimtime="00:00:42.07" resultid="5494" heatid="4866" lane="3" entrytime="00:00:42.87" />
                <RESULT eventid="1175" points="232" reactiontime="0" swimtime="00:00:46.42" resultid="5495" heatid="4897" lane="3" entrytime="00:00:49.76" />
                <RESULT eventid="1267" points="259" reactiontime="0" swimtime="00:00:35.93" resultid="5496" heatid="4927" lane="3" entrytime="00:00:36.82" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Thalles" lastname="Corassari Boas" birthdate="2014-03-10" gender="M" nation="BRA" license="392159" swrid="5466536" athleteid="4833" externalid="392159">
              <RESULTS>
                <RESULT eventid="1090" points="61" reactiontime="0" swimtime="00:00:56.44" resultid="5528" heatid="4860" lane="3" />
                <RESULT eventid="1258" points="55" reactiontime="0" swimtime="00:00:52.92" resultid="5529" heatid="4917" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adan" lastname="Miguel Urdaneta" birthdate="2006-06-08" gender="M" nation="BRA" license="371315" swrid="5603875" athleteid="4794" externalid="371315">
              <RESULTS>
                <RESULT eventid="1135" points="313" reactiontime="0" swimtime="00:01:06.02" resultid="5508" heatid="4884" lane="2" entrytime="00:01:08.94" />
                <RESULT eventid="1275" points="274" reactiontime="0" swimtime="00:00:31.01" resultid="5509" heatid="4931" lane="5" entrytime="00:00:30.73" />
                <RESULT eventid="1323" points="313" reactiontime="0" swimtime="00:00:32.00" resultid="5510" heatid="4947" lane="2" entrytime="00:00:33.37" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Augusto Schmidt" birthdate="2009-05-04" gender="M" nation="BRA" license="367087" athleteid="4827" externalid="367087">
              <RESULTS>
                <RESULT eventid="1275" reactiontime="0" status="DNS" swimtime="00:00:00.00" resultid="5503" entrytime="00:00:42.01" />
                <RESULT eventid="1323" reactiontime="0" status="DNS" swimtime="00:00:00.00" resultid="5504" entrytime="00:00:46.15" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Samuel" lastname="Massuda Santos" birthdate="2012-06-09" gender="M" nation="BRA" license="392189" swrid="5603872" athleteid="4846" externalid="392189">
              <RESULTS>
                <RESULT eventid="1096" points="115" reactiontime="0" swimtime="00:00:45.63" resultid="5537" heatid="4863" lane="5" />
                <RESULT eventid="1124" points="110" reactiontime="0" swimtime="00:01:33.52" resultid="5538" heatid="4876" lane="4" />
                <RESULT eventid="1264" points="138" reactiontime="0" swimtime="00:00:38.94" resultid="5539" heatid="4923" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Gomes Ortiz" birthdate="2008-10-11" gender="M" nation="BRA" license="367082" swrid="5603845" athleteid="4786" externalid="367082">
              <RESULTS>
                <RESULT eventid="1183" points="152" reactiontime="0" swimtime="00:00:46.66" resultid="5497" heatid="4899" lane="6" entrytime="00:00:52.01" />
                <RESULT eventid="1275" points="190" reactiontime="0" swimtime="00:00:35.02" resultid="5498" heatid="4930" lane="2" entrytime="00:00:35.97" />
                <RESULT eventid="1323" reactiontime="0" status="DSQ" swimtime="00:00:00.00" resultid="5499" heatid="4945" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Pedro Venâncio" birthdate="2007-11-22" gender="M" nation="BRA" license="371316" swrid="5603891" athleteid="4810" externalid="371316">
              <RESULTS>
                <RESULT eventid="1275" points="260" reactiontime="0" swimtime="00:00:31.55" resultid="5520" heatid="4930" lane="6" entrytime="00:00:34.72" />
                <RESULT eventid="1323" points="206" reactiontime="0" swimtime="00:00:36.77" resultid="5521" heatid="4946" lane="4" entrytime="00:00:38.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Lucas De Miranda Kmita" birthdate="2005-05-04" gender="M" nation="BRA" license="347848" swrid="5603865" athleteid="4790" externalid="347848">
              <RESULTS>
                <RESULT eventid="1135" points="327" reactiontime="0" swimtime="00:01:05.04" resultid="5505" heatid="4884" lane="6" entrytime="00:01:05.43" />
                <RESULT eventid="1275" points="357" reactiontime="0" swimtime="00:00:28.40" resultid="5506" heatid="4932" lane="7" entrytime="00:00:28.27" />
                <RESULT eventid="1323" points="318" reactiontime="0" swimtime="00:00:31.85" resultid="5507" heatid="4947" lane="6" entrytime="00:00:31.74" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Pauloski Murante" birthdate="1997-06-06" gender="M" nation="BRA" license="367086" swrid="5603887" athleteid="4823" externalid="367086">
              <RESULTS>
                <RESULT eventid="1135" points="237" reactiontime="0" swimtime="00:01:12.41" resultid="5500" heatid="4883" lane="5" entrytime="00:01:13.67" />
                <RESULT eventid="1275" points="260" reactiontime="0" swimtime="00:00:31.55" resultid="5501" heatid="4931" lane="3" entrytime="00:00:31.73" />
                <RESULT eventid="1377" points="156" reactiontime="0" swimtime="00:01:42.52" resultid="5502" heatid="4959" lane="4" entrytime="00:01:46.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Ferreira Batista" birthdate="2014-11-26" gender="F" nation="BRA" license="392160" swrid="5515815" athleteid="4836" externalid="392160">
              <RESULTS>
                <RESULT eventid="1087" reactiontime="0" status="DNS" swimtime="00:00:00.00" resultid="5530" />
                <RESULT eventid="1255" points="48" reactiontime="0" swimtime="00:01:02.88" resultid="5531" heatid="4915" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
