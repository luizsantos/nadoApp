<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.80168">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Maringá" name="Torneio Regional da 2ª Região (Pré-Mirim/Sênior)" course="SCM" deadline="2024-08-13" entrystartdate="2024-08-06" entrytype="INVITATION" hostclub="Universidade Estadual de Maringá" hostclub.url="http://www.uem.br/" number="38313" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/newInterface/eventos/38313" startmethod="2" timing="AUTOMATIC" touchpad="ONESIDE" masters="F" withdrawuntil="2024-08-14" state="PR" nation="BRA" hytek.courseorder="S">
      <AGEDATE value="2024-01-01" type="YEAR" />
      <POOL name="Universidade Estadual de Maringá" lanemin="1" lanemax="6" />
      <FACILITY city="Maringá" name="Universidade Estadual de Maringá" nation="BRA" state="PR" street="M19" street2="Vila Esperança" zip="87020-900" />
      <POINTTABLE pointtableid="3017" name="AQUA Point Scoring" version="2024" />
      <QUALIFY from="2023-08-18" until="2024-08-16" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99252-0598" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99252-0598" street="Avenida do Batel, 1230" street2="Sala 202" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2024-08-17" daytime="09:10" endtime="12:34" number="1" officialmeeting="08:30" teamleadermeeting="09:00" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="1060" daytime="09:10" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1061" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1516" />
                    <RANKING order="2" place="2" resultid="1719" />
                    <RANKING order="3" place="3" resultid="1444" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1699" />
                    <RANKING order="2" place="2" resultid="1757" />
                    <RANKING order="3" place="3" resultid="1847" />
                    <RANKING order="4" place="4" resultid="1440" />
                    <RANKING order="5" place="-1" resultid="1741" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2038" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2039" daytime="09:15" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1063" daytime="09:20" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1064" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1485" />
                    <RANKING order="2" place="2" resultid="1753" />
                    <RANKING order="3" place="3" resultid="1524" />
                    <RANKING order="4" place="4" resultid="1489" />
                    <RANKING order="5" place="5" resultid="1715" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1424" />
                    <RANKING order="2" place="2" resultid="1633" />
                    <RANKING order="3" place="3" resultid="1691" />
                    <RANKING order="4" place="4" resultid="1481" />
                    <RANKING order="5" place="5" resultid="1357" />
                    <RANKING order="6" place="6" resultid="1641" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2040" daytime="09:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2041" daytime="09:25" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1066" daytime="09:30" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1881" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1729" />
                    <RANKING order="2" place="-1" resultid="1331" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1882" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1293" />
                    <RANKING order="2" place="2" resultid="1299" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1883" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1884" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1885" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1320" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1886" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1887" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2042" daytime="09:30" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1070" daytime="09:35" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1888" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1393" />
                    <RANKING order="2" place="2" resultid="1667" />
                    <RANKING order="3" place="3" resultid="1311" />
                    <RANKING order="4" place="-1" resultid="1661" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1889" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1342" />
                    <RANKING order="2" place="2" resultid="1685" />
                    <RANKING order="3" place="3" resultid="1386" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1890" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1891" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1305" />
                    <RANKING order="2" place="2" resultid="1679" />
                    <RANKING order="3" place="3" resultid="1477" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1892" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1277" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1893" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1894" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1820" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2043" daytime="09:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2044" daytime="09:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2045" daytime="09:40" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1077" daytime="09:45" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1078" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1602" />
                    <RANKING order="2" place="2" resultid="1749" />
                    <RANKING order="3" place="3" resultid="1316" />
                    <RANKING order="4" place="4" resultid="1420" />
                    <RANKING order="5" place="5" resultid="1401" />
                    <RANKING order="6" place="6" resultid="1629" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1079" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1619" />
                    <RANKING order="2" place="2" resultid="1416" />
                    <RANKING order="3" place="3" resultid="1700" />
                    <RANKING order="4" place="-1" resultid="1637" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2046" daytime="09:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2047" daytime="09:50" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1080" daytime="09:55" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1081" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1428" />
                    <RANKING order="2" place="2" resultid="1493" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1409" />
                    <RANKING order="2" place="2" resultid="1432" />
                    <RANKING order="3" place="3" resultid="1657" />
                    <RANKING order="4" place="4" resultid="1634" />
                    <RANKING order="5" place="5" resultid="1855" />
                    <RANKING order="6" place="6" resultid="1692" />
                    <RANKING order="7" place="7" resultid="1874" />
                    <RANKING order="8" place="8" resultid="1436" />
                    <RANKING order="9" place="9" resultid="1877" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2048" daytime="09:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2049" daytime="09:55" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1083" daytime="10:00" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1895" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1466" />
                    <RANKING order="2" place="2" resultid="1397" />
                    <RANKING order="3" place="3" resultid="1405" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1896" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1651" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1897" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1898" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1373" />
                    <RANKING order="2" place="2" resultid="1283" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1899" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1289" />
                    <RANKING order="2" place="2" resultid="1361" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1900" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1826" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1901" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1575" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2050" daytime="10:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2051" daytime="10:00" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1091" daytime="10:05" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1092" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1390" />
                    <RANKING order="2" place="2" resultid="1674" />
                    <RANKING order="3" place="3" resultid="1614" />
                    <RANKING order="4" place="4" resultid="1463" />
                    <RANKING order="5" place="-1" resultid="1623" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1093" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1504" />
                    <RANKING order="2" place="2" resultid="1326" />
                    <RANKING order="3" place="3" resultid="1865" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1382" />
                    <RANKING order="2" place="2" resultid="1836" />
                    <RANKING order="3" place="3" resultid="1816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1095" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1378" />
                    <RANKING order="2" place="2" resultid="1350" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1096" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1831" />
                    <RANKING order="2" place="-1" resultid="1579" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1097" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1842" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1821" />
                    <RANKING order="2" place="2" resultid="1338" />
                    <RANKING order="3" place="3" resultid="1555" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2052" daytime="10:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2053" daytime="10:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2054" daytime="10:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2055" daytime="10:15" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1099" daytime="10:15" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1100" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1603" />
                    <RANKING order="2" place="2" resultid="1517" />
                    <RANKING order="3" place="3" resultid="1703" />
                    <RANKING order="4" place="4" resultid="1750" />
                    <RANKING order="5" place="5" resultid="1707" />
                    <RANKING order="6" place="6" resultid="1317" />
                    <RANKING order="7" place="7" resultid="1445" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1101" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1417" />
                    <RANKING order="2" place="2" resultid="1848" />
                    <RANKING order="3" place="3" resultid="1441" />
                    <RANKING order="4" place="-1" resultid="1791" />
                    <RANKING order="5" place="-1" resultid="1742" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2056" daytime="10:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2057" daytime="10:20" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1102" daytime="10:20" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1103" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1486" />
                    <RANKING order="2" place="2" resultid="1525" />
                    <RANKING order="3" place="3" resultid="1716" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1104" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1856" />
                    <RANKING order="2" place="2" resultid="1642" />
                    <RANKING order="3" place="3" resultid="1358" />
                    <RANKING order="4" place="4" resultid="1482" />
                    <RANKING order="5" place="5" resultid="1804" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2058" daytime="10:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2059" daytime="10:25" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1105" daytime="10:25" gender="F" number="11" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1902" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1731" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1903" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1904" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1905" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1906" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1608" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1907" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1908" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2060" daytime="10:25" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1109" daytime="10:50" gender="M" number="12" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1909" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1613" />
                    <RANKING order="2" place="2" resultid="1673" />
                    <RANKING order="3" place="3" resultid="1668" />
                    <RANKING order="4" place="-1" resultid="1662" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1910" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2144" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1911" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2146" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1912" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2145" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1913" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1914" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1915" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2061" daytime="10:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2062" daytime="11:10" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1114" daytime="11:40" gender="F" number="13" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1115" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1518" />
                    <RANKING order="2" place="2" resultid="1708" />
                    <RANKING order="3" place="3" resultid="1720" />
                    <RANKING order="4" place="4" resultid="1402" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1116" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1758" />
                    <RANKING order="2" place="-1" resultid="1792" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2063" daytime="11:40" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1117" daytime="11:45" gender="M" number="14" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1118" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1754" />
                    <RANKING order="2" place="2" resultid="1429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1119" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1433" />
                    <RANKING order="2" place="2" resultid="1426" />
                    <RANKING order="3" place="3" resultid="1410" />
                    <RANKING order="4" place="4" resultid="1635" />
                    <RANKING order="5" place="5" resultid="1693" />
                    <RANKING order="6" place="6" resultid="1658" />
                    <RANKING order="7" place="7" resultid="1805" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2064" daytime="11:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2065" daytime="11:45" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1120" daytime="11:50" gender="F" number="15" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1916" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1332" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1917" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1859" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1918" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1919" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1920" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1607" />
                    <RANKING order="2" place="2" resultid="1362" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1921" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1922" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1808" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2066" daytime="11:50" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1126" daytime="11:55" gender="M" number="16" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1923" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1924" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1925" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1926" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1927" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1278" />
                    <RANKING order="2" place="2" resultid="1832" />
                    <RANKING order="3" place="-1" resultid="1580" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1928" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1929" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2067" daytime="11:55" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1128" daytime="11:55" gender="F" number="17" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1129" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1721" />
                    <RANKING order="2" place="2" resultid="1704" />
                    <RANKING order="3" place="3" resultid="1446" />
                    <RANKING order="4" place="4" resultid="1421" />
                    <RANKING order="5" place="5" resultid="1630" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1130" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1442" />
                    <RANKING order="2" place="2" resultid="1759" />
                    <RANKING order="3" place="-1" resultid="1620" />
                    <RANKING order="4" place="-1" resultid="1638" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2068" daytime="11:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2069" daytime="12:00" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1131" daytime="12:05" gender="M" number="18" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1132" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1487" />
                    <RANKING order="2" place="2" resultid="1494" />
                    <RANKING order="3" place="3" resultid="1490" />
                    <RANKING order="4" place="4" resultid="1526" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1133" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1425" />
                    <RANKING order="2" place="2" resultid="1359" />
                    <RANKING order="3" place="-1" resultid="1437" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2070" daytime="12:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2071" daytime="12:10" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1134" daytime="12:15" gender="F" number="19" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1930" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1730" />
                    <RANKING order="2" place="-1" resultid="1398" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1931" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1455" />
                    <RANKING order="2" place="2" resultid="1300" />
                    <RANKING order="3" place="3" resultid="1294" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1932" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1370" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1933" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1285" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1934" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1322" />
                    <RANKING order="2" place="2" resultid="1291" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1935" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1936" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2072" daytime="12:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2073" daytime="12:20" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1140" daytime="12:20" gender="M" number="20" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1937" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1669" />
                    <RANKING order="2" place="2" resultid="1354" />
                    <RANKING order="3" place="-1" resultid="1663" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1938" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1939" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1646" />
                    <RANKING order="2" place="2" resultid="1413" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1940" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1469" />
                    <RANKING order="2" place="2" resultid="1681" />
                    <RANKING order="3" place="-1" resultid="1306" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1941" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1942" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1943" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2074" daytime="12:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2075" daytime="12:25" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1144" daytime="12:30" gender="F" number="21" order="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1145" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1604" />
                    <RANKING order="2" place="2" resultid="1751" />
                    <RANKING order="3" place="3" resultid="1318" />
                    <RANKING order="4" place="4" resultid="1709" />
                    <RANKING order="5" place="5" resultid="1705" />
                    <RANKING order="6" place="6" resultid="1403" />
                    <RANKING order="7" place="7" resultid="1631" />
                    <RANKING order="8" place="8" resultid="1727" />
                    <RANKING order="9" place="9" resultid="1422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1146" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1621" />
                    <RANKING order="2" place="2" resultid="1418" />
                    <RANKING order="3" place="3" resultid="1849" />
                    <RANKING order="4" place="4" resultid="1701" />
                    <RANKING order="5" place="5" resultid="1793" />
                    <RANKING order="6" place="-1" resultid="1639" />
                    <RANKING order="7" place="-1" resultid="1743" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2076" daytime="12:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2077" daytime="12:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2078" daytime="12:30" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1147" daytime="12:35" gender="M" number="22" order="23" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1148" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1755" />
                    <RANKING order="2" place="2" resultid="1495" />
                    <RANKING order="3" place="3" resultid="1491" />
                    <RANKING order="4" place="4" resultid="1430" />
                    <RANKING order="5" place="5" resultid="1717" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1149" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1434" />
                    <RANKING order="2" place="2" resultid="1411" />
                    <RANKING order="3" place="3" resultid="1659" />
                    <RANKING order="4" place="4" resultid="1857" />
                    <RANKING order="5" place="5" resultid="1438" />
                    <RANKING order="6" place="6" resultid="1483" />
                    <RANKING order="7" place="7" resultid="1643" />
                    <RANKING order="8" place="8" resultid="1875" />
                    <RANKING order="9" place="9" resultid="1878" />
                    <RANKING order="10" place="10" resultid="1806" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2079" daytime="12:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2080" daytime="12:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2081" daytime="12:35" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1150" daytime="12:40" gender="F" number="23" order="24" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1944" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1945" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1452" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1946" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1947" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1284" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1948" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1321" />
                    <RANKING order="2" place="-1" resultid="1290" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1949" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1827" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1950" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1576" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2082" daytime="12:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2083" daytime="12:40" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1157" daytime="12:45" gender="M" number="24" order="25" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1951" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1394" />
                    <RANKING order="2" place="2" resultid="1312" />
                    <RANKING order="3" place="3" resultid="1812" />
                    <RANKING order="4" place="-1" resultid="1870" />
                    <RANKING order="5" place="-1" resultid="1624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1952" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1687" />
                    <RANKING order="2" place="2" resultid="1866" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1953" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1837" />
                    <RANKING order="2" place="2" resultid="1414" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1954" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1379" />
                    <RANKING order="2" place="2" resultid="1478" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1955" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1279" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1956" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1843" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1957" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1339" />
                    <RANKING order="2" place="2" resultid="1822" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2084" daytime="12:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2085" daytime="12:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2086" daytime="12:45" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-08-17" daytime="15:40" endtime="18:06" number="2" officialmeeting="15:00" teamleadermeeting="15:30" warmupfrom="14:30" warmupuntil="15:30">
          <EVENTS>
            <EVENT eventid="1165" daytime="15:40" gender="F" number="25" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1166" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1583" />
                    <RANKING order="2" place="2" resultid="1797" />
                    <RANKING order="3" place="-1" resultid="1597" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2087" daytime="15:40" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1167" daytime="15:40" gender="M" number="26" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2028" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1776" />
                    <RANKING order="2" place="2" resultid="1566" />
                    <RANKING order="3" place="3" resultid="1592" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2088" daytime="15:40" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1169" daytime="15:45" gender="F" number="27" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1170" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1588" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1171" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1695" />
                    <RANKING order="2" place="2" resultid="1851" />
                    <RANKING order="3" place="-1" resultid="1711" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2089" daytime="15:45" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1172" daytime="15:45" gender="M" number="28" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1173" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1528" />
                    <RANKING order="2" place="2" resultid="1473" />
                    <RANKING order="3" place="3" resultid="1512" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1174" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1520" />
                    <RANKING order="2" place="2" resultid="1459" />
                    <RANKING order="3" place="3" resultid="1764" />
                    <RANKING order="4" place="4" resultid="1508" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2090" daytime="15:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2091" daytime="15:50" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1175" daytime="15:55" gender="F" number="29" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1958" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1406" />
                    <RANKING order="2" place="2" resultid="1732" />
                    <RANKING order="3" place="-1" resultid="1333" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1959" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1295" />
                    <RANKING order="2" place="2" resultid="1456" />
                    <RANKING order="3" place="3" resultid="1301" />
                    <RANKING order="4" place="4" resultid="1653" />
                    <RANKING order="5" place="5" resultid="1860" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1960" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1961" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1375" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1962" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1609" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1963" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1964" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2092" daytime="15:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2093" daytime="16:00" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1180" daytime="16:10" gender="M" number="30" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1965" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1395" />
                    <RANKING order="2" place="2" resultid="1675" />
                    <RANKING order="3" place="3" resultid="1615" />
                    <RANKING order="4" place="4" resultid="1670" />
                    <RANKING order="5" place="5" resultid="1768" />
                    <RANKING order="6" place="6" resultid="1625" />
                    <RANKING order="7" place="-1" resultid="1664" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1966" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1343" />
                    <RANKING order="2" place="2" resultid="1688" />
                    <RANKING order="3" place="3" resultid="1505" />
                    <RANKING order="4" place="4" resultid="1867" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1967" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1647" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1968" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1351" />
                    <RANKING order="2" place="2" resultid="1479" />
                    <RANKING order="3" place="3" resultid="1682" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1969" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1970" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1971" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1880" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2094" daytime="16:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2095" daytime="16:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2096" daytime="16:20" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1186" daytime="16:30" gender="F" number="31" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2029" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1584" />
                    <RANKING order="2" place="2" resultid="1798" />
                    <RANKING order="3" place="3" resultid="1780" />
                    <RANKING order="4" place="4" resultid="1784" />
                    <RANKING order="5" place="-1" resultid="1598" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2097" daytime="16:30" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1188" daytime="16:30" gender="M" number="32" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2030" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1593" />
                    <RANKING order="2" place="2" resultid="1777" />
                    <RANKING order="3" place="3" resultid="1567" />
                    <RANKING order="4" place="-1" resultid="1788" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2098" daytime="16:30" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1190" daytime="16:30" gender="F" number="33" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1191" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1547" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1192" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1696" />
                    <RANKING order="2" place="2" resultid="1551" />
                    <RANKING order="3" place="3" resultid="1540" />
                    <RANKING order="4" place="4" resultid="1558" />
                    <RANKING order="5" place="5" resultid="1852" />
                    <RANKING order="6" place="-1" resultid="1745" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2099" daytime="16:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2100" daytime="16:35" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1193" daytime="16:35" gender="M" number="34" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1194" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1529" />
                    <RANKING order="2" place="2" resultid="1735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1195" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1460" />
                    <RANKING order="2" place="2" resultid="1509" />
                    <RANKING order="3" place="3" resultid="1772" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2101" daytime="16:35" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1196" daytime="16:40" gender="F" number="35" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1972" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1501" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1973" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1453" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1974" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1975" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1365" />
                    <RANKING order="2" place="2" resultid="1286" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1976" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1323" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1977" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1828" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1978" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2102" daytime="16:40" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1202" daytime="16:45" gender="M" number="36" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1979" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1355" />
                    <RANKING order="2" place="2" resultid="1313" />
                    <RANKING order="3" place="3" resultid="1626" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1980" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1689" />
                    <RANKING order="2" place="2" resultid="1387" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1981" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1348" />
                    <RANKING order="2" place="2" resultid="1838" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1982" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1307" />
                    <RANKING order="2" place="2" resultid="1352" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1983" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1280" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1984" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1844" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1985" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2103" daytime="16:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2104" daytime="16:45" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1209" daytime="17:05" gender="F" number="37" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2031" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1585" />
                    <RANKING order="2" place="2" resultid="1785" />
                    <RANKING order="3" place="3" resultid="1781" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2105" daytime="17:05" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1211" daytime="17:05" gender="M" number="38" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2032" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1568" />
                    <RANKING order="2" place="2" resultid="1594" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2106" daytime="17:05" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1213" daytime="17:10" gender="F" number="39" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1214" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1737" />
                    <RANKING order="2" place="2" resultid="1548" />
                    <RANKING order="3" place="3" resultid="1571" />
                    <RANKING order="4" place="4" resultid="1532" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1215" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1552" />
                    <RANKING order="2" place="2" resultid="1697" />
                    <RANKING order="3" place="3" resultid="1448" />
                    <RANKING order="4" place="4" resultid="2139" />
                    <RANKING order="5" place="5" resultid="1544" />
                    <RANKING order="6" place="-1" resultid="1712" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2107" daytime="17:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2108" daytime="17:10" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1216" daytime="17:15" gender="M" number="40" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1217" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1723" />
                    <RANKING order="2" place="2" resultid="1513" />
                    <RANKING order="3" place="3" resultid="1562" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1218" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1521" />
                    <RANKING order="2" place="2" resultid="1536" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2109" daytime="17:15" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1219" daytime="17:15" gender="F" number="41" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1986" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1334" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1987" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1302" />
                    <RANKING order="2" place="2" resultid="1296" />
                    <RANKING order="3" place="3" resultid="1861" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1988" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1371" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1989" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1376" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1990" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1610" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1991" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1992" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2110" daytime="17:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2111" daytime="17:20" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1225" daytime="17:20" gender="M" number="42" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1993" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1671" />
                    <RANKING order="2" place="2" resultid="1464" />
                    <RANKING order="3" place="3" resultid="1871" />
                    <RANKING order="4" place="4" resultid="1769" />
                    <RANKING order="5" place="5" resultid="1813" />
                    <RANKING order="6" place="-1" resultid="1616" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1994" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1327" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1995" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1383" />
                    <RANKING order="2" place="2" resultid="1648" />
                    <RANKING order="3" place="3" resultid="1839" />
                    <RANKING order="4" place="4" resultid="1817" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1996" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1308" />
                    <RANKING order="2" place="2" resultid="1470" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1997" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1998" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1999" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1823" />
                    <RANKING order="2" place="2" resultid="1497" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2112" daytime="17:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2113" daytime="17:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2114" daytime="17:25" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1231" daytime="17:25" gender="F" number="43" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2033" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1586" />
                    <RANKING order="2" place="2" resultid="1799" />
                    <RANKING order="3" place="3" resultid="1786" />
                    <RANKING order="4" place="4" resultid="1782" />
                    <RANKING order="5" place="-1" resultid="1599" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2115" daytime="17:25" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1233" daytime="17:30" gender="M" number="44" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2034" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1778" />
                    <RANKING order="2" place="2" resultid="1595" />
                    <RANKING order="3" place="3" resultid="1569" />
                    <RANKING order="4" place="-1" resultid="1789" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2116" daytime="17:30" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1235" daytime="17:30" gender="F" number="45" order="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1236" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1589" />
                    <RANKING order="2" place="2" resultid="1738" />
                    <RANKING order="3" place="3" resultid="1572" />
                    <RANKING order="4" place="4" resultid="1533" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1237" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1449" />
                    <RANKING order="2" place="2" resultid="1761" />
                    <RANKING order="3" place="3" resultid="1559" />
                    <RANKING order="4" place="4" resultid="1541" />
                    <RANKING order="5" place="-1" resultid="1746" />
                    <RANKING order="6" place="-1" resultid="1853" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2117" daytime="17:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2118" daytime="17:35" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1238" daytime="17:35" gender="M" number="46" order="23" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1239" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1530" />
                    <RANKING order="2" place="2" resultid="1474" />
                    <RANKING order="3" place="3" resultid="1563" />
                    <RANKING order="4" place="4" resultid="1724" />
                    <RANKING order="5" place="5" resultid="1514" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1240" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1461" />
                    <RANKING order="2" place="2" resultid="1773" />
                    <RANKING order="3" place="3" resultid="1537" />
                    <RANKING order="4" place="4" resultid="1765" />
                    <RANKING order="5" place="5" resultid="1510" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2119" daytime="17:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2120" daytime="17:40" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1241" daytime="17:40" gender="F" number="47" order="24" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2000" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1467" />
                    <RANKING order="2" place="2" resultid="1407" />
                    <RANKING order="3" place="3" resultid="1733" />
                    <RANKING order="4" place="4" resultid="1502" />
                    <RANKING order="5" place="-1" resultid="1399" />
                    <RANKING order="6" place="-1" resultid="1335" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2001" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1654" />
                    <RANKING order="2" place="2" resultid="1862" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2002" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1368" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2003" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1287" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2004" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1324" />
                    <RANKING order="2" place="2" resultid="1611" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2005" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="2006" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1809" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2121" daytime="17:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2122" daytime="17:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2123" daytime="17:50" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1248" daytime="17:50" gender="M" number="48" order="25" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2007" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1391" />
                    <RANKING order="2" place="2" resultid="1676" />
                    <RANKING order="3" place="-1" resultid="1617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2008" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1388" />
                    <RANKING order="2" place="2" resultid="1506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2009" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1384" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2010" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1683" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2011" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1281" />
                    <RANKING order="2" place="2" resultid="1833" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2012" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="2013" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2124" daytime="17:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2125" daytime="17:55" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1254" daytime="18:00" gender="F" number="49" order="26" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1255" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1549" />
                    <RANKING order="2" place="2" resultid="1590" />
                    <RANKING order="3" place="3" resultid="1739" />
                    <RANKING order="4" place="4" resultid="1573" />
                    <RANKING order="5" place="5" resultid="1534" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1256" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1553" />
                    <RANKING order="2" place="2" resultid="1801" />
                    <RANKING order="3" place="3" resultid="1450" />
                    <RANKING order="4" place="4" resultid="1762" />
                    <RANKING order="5" place="5" resultid="1542" />
                    <RANKING order="6" place="6" resultid="1545" />
                    <RANKING order="7" place="-1" resultid="1560" />
                    <RANKING order="8" place="-1" resultid="1713" />
                    <RANKING order="9" place="-1" resultid="1747" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2126" daytime="18:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2127" daytime="18:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2128" daytime="18:00" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1257" daytime="18:05" gender="M" number="50" order="27" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1258" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1725" />
                    <RANKING order="2" place="2" resultid="1475" />
                    <RANKING order="3" place="3" resultid="1564" />
                    <RANKING order="4" place="-1" resultid="1795" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1259" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1522" />
                    <RANKING order="2" place="2" resultid="1538" />
                    <RANKING order="3" place="3" resultid="1774" />
                    <RANKING order="4" place="4" resultid="1766" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2129" daytime="18:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2130" daytime="18:05" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1260" daytime="18:10" gender="F" number="51" order="28" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2014" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="2015" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1457" />
                    <RANKING order="2" place="2" resultid="1303" />
                    <RANKING order="3" place="3" resultid="1297" />
                    <RANKING order="4" place="4" resultid="1655" />
                    <RANKING order="5" place="5" resultid="1863" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2016" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="2017" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="2018" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1363" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2019" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1829" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2020" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1810" />
                    <RANKING order="2" place="2" resultid="1577" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2131" daytime="18:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2132" daytime="18:10" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1265" daytime="18:15" gender="M" number="52" order="29" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2021" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1665" />
                    <RANKING order="2" place="2" resultid="1677" />
                    <RANKING order="3" place="3" resultid="1314" />
                    <RANKING order="4" place="4" resultid="1627" />
                    <RANKING order="5" place="5" resultid="1872" />
                    <RANKING order="6" place="6" resultid="1770" />
                    <RANKING order="7" place="7" resultid="1814" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2022" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1328" />
                    <RANKING order="2" place="2" resultid="1868" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2023" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1840" />
                    <RANKING order="2" place="2" resultid="1649" />
                    <RANKING order="3" place="3" resultid="1818" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2024" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1345" />
                    <RANKING order="2" place="2" resultid="1309" />
                    <RANKING order="3" place="3" resultid="1471" />
                    <RANKING order="4" place="-1" resultid="1380" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2025" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1834" />
                    <RANKING order="2" place="2" resultid="1581" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2026" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1845" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2027" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1340" />
                    <RANKING order="2" place="2" resultid="1824" />
                    <RANKING order="3" place="3" resultid="1556" />
                    <RANKING order="4" place="4" resultid="1498" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2133" daytime="18:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2134" daytime="18:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2135" daytime="18:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2136" daytime="18:20" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="1035" nation="BRA" region="PR" clubid="1802" swrid="93778" name="Fundação De Esportes De Campo Mourão" shortname="Fecam">
          <ATHLETES>
            <ATHLETE firstname="Beatriz" lastname="Ferreira Batista" birthdate="2014-11-26" gender="F" nation="BRA" license="392160" swrid="5515815" athleteid="1850" externalid="392160">
              <RESULTS>
                <RESULT eventid="1169" points="95" swimtime="00:01:50.00" resultid="1851" heatid="2089" lane="5" />
                <RESULT eventid="1190" points="27" swimtime="00:01:20.79" resultid="1852" heatid="2099" lane="2" />
                <RESULT eventid="1235" status="DNS" swimtime="00:00:00.00" resultid="1853" heatid="2117" lane="2" />
                <RESULT eventid="1213" points="94" swimtime="00:00:55.39" resultid="2139" heatid="2107" lane="5" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Giroldo Santos" birthdate="2011-05-16" gender="M" nation="BRA" license="399602" athleteid="1869" externalid="399602">
              <RESULTS>
                <RESULT eventid="1157" status="DSQ" swimtime="00:00:49.36" resultid="1870" heatid="2085" lane="1" />
                <RESULT eventid="1225" points="155" swimtime="00:00:40.47" resultid="1871" heatid="2112" lane="4" />
                <RESULT eventid="1265" points="201" swimtime="00:00:34.40" resultid="1872" heatid="2134" lane="4" entrytime="00:00:35.31" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Keirrison" lastname="Leite Silva" birthdate="2011-08-02" gender="M" nation="BRA" license="392161" swrid="5603864" athleteid="1811" externalid="392161">
              <RESULTS>
                <RESULT eventid="1157" points="98" swimtime="00:00:53.97" resultid="1812" heatid="2085" lane="5" />
                <RESULT eventid="1225" points="64" swimtime="00:00:54.23" resultid="1813" heatid="2113" lane="1" />
                <RESULT eventid="1265" points="106" swimtime="00:00:42.57" resultid="1814" heatid="2133" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Samuel" lastname="Massuda Santos" birthdate="2012-06-09" gender="M" nation="BRA" license="392189" swrid="5603872" athleteid="1854" externalid="392189">
              <RESULTS>
                <RESULT eventid="1080" points="162" swimtime="00:01:41.32" resultid="1855" heatid="2049" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="165" swimtime="00:00:40.28" resultid="1856" heatid="2059" lane="2" />
                <RESULT eventid="1147" points="209" swimtime="00:00:33.95" resultid="1857" heatid="2081" lane="2" entrytime="00:00:33.62" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Gabrieli Oliveira" birthdate="2010-09-23" gender="F" nation="BRA" license="403428" swrid="5676288" athleteid="1858" externalid="403428">
              <RESULTS>
                <RESULT eventid="1120" points="196" swimtime="00:00:43.45" resultid="1859" heatid="2066" lane="5" entrytime="00:00:44.54" entrycourse="SCM" />
                <RESULT eventid="1175" points="206" swimtime="00:06:31.06" resultid="1860" heatid="2092" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.03" />
                    <SPLIT distance="100" swimtime="00:01:24.67" />
                    <SPLIT distance="150" swimtime="00:02:15.48" />
                    <SPLIT distance="200" swimtime="00:03:04.89" />
                    <SPLIT distance="250" swimtime="00:03:56.06" />
                    <SPLIT distance="300" swimtime="00:04:48.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="172" swimtime="00:00:43.78" resultid="1861" heatid="2110" lane="4" />
                <RESULT eventid="1241" points="193" swimtime="00:01:34.98" resultid="1862" heatid="2122" lane="2" entrytime="00:01:34.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1260" points="271" swimtime="00:00:35.42" resultid="1863" heatid="2132" lane="6" entrytime="00:00:35.41" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Felipe Damha" birthdate="1987-01-02" gender="M" nation="BRA" license="053982" athleteid="1879" externalid="053982">
              <RESULTS>
                <RESULT eventid="1180" points="304" swimtime="00:05:15.57" resultid="1880" heatid="2095" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                    <SPLIT distance="100" swimtime="00:01:12.75" />
                    <SPLIT distance="150" swimtime="00:01:51.13" />
                    <SPLIT distance="200" swimtime="00:02:30.63" />
                    <SPLIT distance="250" swimtime="00:03:10.55" />
                    <SPLIT distance="300" swimtime="00:03:52.18" />
                    <SPLIT distance="350" swimtime="00:04:34.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kenzo" lastname="Kimura" birthdate="2010-04-23" gender="M" nation="BRA" license="403429" swrid="5676289" athleteid="1864" externalid="403429">
              <RESULTS>
                <RESULT eventid="1091" points="176" swimtime="00:01:19.95" resultid="1865" heatid="2052" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="149" swimtime="00:00:46.96" resultid="1866" heatid="2085" lane="2" />
                <RESULT eventid="1180" points="165" swimtime="00:06:26.41" resultid="1867" heatid="2094" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.53" />
                    <SPLIT distance="100" swimtime="00:01:25.63" />
                    <SPLIT distance="150" swimtime="00:02:15.13" />
                    <SPLIT distance="200" swimtime="00:03:04.79" />
                    <SPLIT distance="250" swimtime="00:03:56.88" />
                    <SPLIT distance="300" swimtime="00:04:48.53" />
                    <SPLIT distance="350" swimtime="00:05:38.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="171" swimtime="00:00:36.28" resultid="1868" heatid="2133" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique De Oliveira" birthdate="2009-07-28" gender="M" nation="BRA" license="414505" athleteid="1815" externalid="414505">
              <RESULTS>
                <RESULT eventid="1091" points="266" swimtime="00:01:09.71" resultid="1816" heatid="2054" lane="4" entrytime="00:01:07.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="337" swimtime="00:00:31.24" resultid="1817" heatid="2114" lane="2" entrytime="00:00:32.62" entrycourse="SCM" />
                <RESULT eventid="1265" points="308" swimtime="00:00:29.82" resultid="1818" heatid="2135" lane="2" entrytime="00:00:29.25" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Eduardo Schork Filho" birthdate="2012-12-28" gender="M" nation="BRA" license="413906" athleteid="1873" externalid="413906">
              <RESULTS>
                <RESULT eventid="1080" points="102" swimtime="00:01:58.13" resultid="1874" heatid="2048" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="107" swimtime="00:00:42.42" resultid="1875" heatid="2079" lane="3" entrytime="00:00:44.28" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Batinga Ponchielli" birthdate="2007-01-18" gender="M" nation="BRA" license="378461" swrid="5251143" athleteid="1830" externalid="378461">
              <RESULTS>
                <RESULT eventid="1091" points="279" swimtime="00:01:08.56" resultid="1831" heatid="2053" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1126" points="243" swimtime="00:00:35.39" resultid="1832" heatid="2067" lane="3" entrytime="00:00:33.52" entrycourse="SCM" />
                <RESULT eventid="1248" points="219" swimtime="00:01:20.14" resultid="1833" heatid="2125" lane="1" entrytime="00:01:18.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="277" swimtime="00:00:30.92" resultid="1834" heatid="2135" lane="1" entrytime="00:00:30.02" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Franca Rebollo" birthdate="2012-09-26" gender="M" nation="BRA" license="385780" swrid="5538081" athleteid="1803" externalid="385780">
              <RESULTS>
                <RESULT eventid="1102" points="83" swimtime="00:00:50.61" resultid="1804" heatid="2058" lane="3" />
                <RESULT eventid="1117" points="73" swimtime="00:01:54.21" resultid="1805" heatid="2065" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="95" swimtime="00:00:44.05" resultid="1806" heatid="2080" lane="6" entrytime="00:00:43.18" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Ferreira Batista" birthdate="2012-03-29" gender="F" nation="BRA" license="385779" swrid="5532525" athleteid="1846" externalid="385779">
              <RESULTS>
                <RESULT eventid="1060" points="229" swimtime="00:03:00.25" resultid="1847" heatid="2038" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.70" />
                    <SPLIT distance="100" swimtime="00:01:28.95" />
                    <SPLIT distance="150" swimtime="00:02:15.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="234" swimtime="00:00:40.97" resultid="1848" heatid="2057" lane="6" entrytime="00:00:44.39" entrycourse="SCM" />
                <RESULT eventid="1144" points="261" swimtime="00:00:35.85" resultid="1849" heatid="2077" lane="2" entrytime="00:00:38.12" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Franco Santos" birthdate="2002-01-03" gender="M" nation="BRA" license="290441" swrid="5546064" athleteid="1819" externalid="290441">
              <RESULTS>
                <RESULT eventid="1070" points="384" swimtime="00:02:30.82" resultid="1820" heatid="2043" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                    <SPLIT distance="100" swimtime="00:01:08.60" />
                    <SPLIT distance="150" swimtime="00:01:55.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1091" points="454" swimtime="00:00:58.34" resultid="1821" heatid="2055" lane="3" entrytime="00:00:56.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="463" swimtime="00:00:32.25" resultid="1822" heatid="2084" lane="3" />
                <RESULT eventid="1225" points="501" swimtime="00:00:27.37" resultid="1823" heatid="2114" lane="3" entrytime="00:00:27.76" entrycourse="SCM" />
                <RESULT eventid="1265" points="499" swimtime="00:00:25.41" resultid="1824" heatid="2136" lane="3" entrytime="00:00:25.79" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Stipp Silva" birthdate="2009-12-02" gender="M" nation="BRA" license="378462" swrid="5603918" athleteid="1835" externalid="378462">
              <RESULTS>
                <RESULT eventid="1091" points="398" swimtime="00:01:00.95" resultid="1836" heatid="2055" lane="2" entrytime="00:01:02.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="316" swimtime="00:00:36.60" resultid="1837" heatid="2086" lane="6" entrytime="00:00:39.01" entrycourse="SCM" />
                <RESULT eventid="1202" points="308" swimtime="00:01:21.83" resultid="1838" heatid="2103" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="358" swimtime="00:00:30.63" resultid="1839" heatid="2113" lane="6" />
                <RESULT eventid="1265" points="421" swimtime="00:00:26.88" resultid="1840" heatid="2136" lane="5" entrytime="00:00:27.52" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Gomes De Souza" birthdate="2006-01-30" gender="F" nation="BRA" license="308464" swrid="5603844" athleteid="1825" externalid="308464">
              <RESULTS>
                <RESULT eventid="1083" points="233" swimtime="00:01:21.64" resultid="1826" heatid="2050" lane="4" entrytime="00:01:19.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1150" points="283" swimtime="00:00:43.19" resultid="1827" heatid="2083" lane="4" entrytime="00:00:43.86" entrycourse="SCM" />
                <RESULT eventid="1196" points="204" swimtime="00:01:45.92" resultid="1828" heatid="2102" lane="6" entrytime="00:01:41.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1260" points="294" swimtime="00:00:34.47" resultid="1829" heatid="2132" lane="1" entrytime="00:00:33.91" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaue" lastname="Guilherme Chagas" birthdate="2005-06-29" gender="M" nation="BRA" license="378464" swrid="5603851" athleteid="1841" externalid="378464">
              <RESULTS>
                <RESULT eventid="1091" points="368" swimtime="00:01:02.52" resultid="1842" heatid="2055" lane="1" entrytime="00:01:04.01" entrycourse="SCM" />
                <RESULT eventid="1157" points="259" swimtime="00:00:39.14" resultid="1843" heatid="2085" lane="6" />
                <RESULT eventid="1202" points="256" swimtime="00:01:26.99" resultid="1844" heatid="2103" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="348" swimtime="00:00:28.65" resultid="1845" heatid="2135" lane="3" entrytime="00:00:29.14" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henry" lastname="Sadao Da Silva" birthdate="2012-10-02" gender="M" nation="BRA" license="413907" athleteid="1876" externalid="413907">
              <RESULTS>
                <RESULT eventid="1080" points="70" swimtime="00:02:13.80" resultid="1877" heatid="2048" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="99" swimtime="00:00:43.55" resultid="1878" heatid="2079" lane="4" entrytime="00:00:46.84" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduarda" lastname="Daleffe Pepino" birthdate="2000-07-09" gender="F" nation="BRA" license="185817" athleteid="1807" externalid="185817">
              <RESULTS>
                <RESULT eventid="1120" points="364" swimtime="00:00:35.34" resultid="1808" heatid="2066" lane="6" />
                <RESULT eventid="1241" points="296" swimtime="00:01:22.33" resultid="1809" heatid="2121" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1260" points="380" swimtime="00:00:31.65" resultid="1810" heatid="2131" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15981" nation="BRA" region="PR" clubid="1275" swrid="93783" name="Quinto Nado" shortname="5º Nado">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Fernanda Romero" birthdate="2007-04-18" gender="F" nation="BRA" license="404750" swrid="4828153" athleteid="1319" externalid="404750">
              <RESULTS>
                <RESULT eventid="1066" points="496" swimtime="00:02:33.94" resultid="1320" heatid="2042" lane="3" entrytime="00:02:34.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                    <SPLIT distance="100" swimtime="00:01:14.26" />
                    <SPLIT distance="150" swimtime="00:01:58.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1150" points="504" swimtime="00:00:35.64" resultid="1321" heatid="2083" lane="5" />
                <RESULT eventid="1134" points="459" swimtime="00:01:10.04" resultid="1322" heatid="2073" lane="3" entrytime="00:01:10.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="451" swimtime="00:01:21.30" resultid="1323" heatid="2102" lane="4" entrytime="00:01:19.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1241" points="430" swimtime="00:01:12.68" resultid="1324" heatid="2121" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Betina" lastname="Tramontini Queiroz" birthdate="2007-09-11" gender="F" nation="BRA" license="357155" swrid="5658063" athleteid="1288" externalid="357155" level="VIBE">
              <RESULTS>
                <RESULT eventid="1083" points="430" swimtime="00:01:06.57" resultid="1289" heatid="2051" lane="3" entrytime="00:01:02.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1150" status="DNS" swimtime="00:00:00.00" resultid="1290" heatid="2082" lane="2" />
                <RESULT eventid="1134" points="310" swimtime="00:01:19.79" resultid="1291" heatid="2073" lane="2" entrytime="00:01:17.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="Sorace Spironelli" birthdate="2008-05-14" gender="M" nation="BRA" license="371318" swrid="5622308" athleteid="1304" externalid="371318">
              <RESULTS>
                <RESULT eventid="1070" points="377" swimtime="00:02:31.75" resultid="1305" heatid="2043" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                    <SPLIT distance="100" swimtime="00:01:11.81" />
                    <SPLIT distance="150" swimtime="00:01:55.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" status="DSQ" swimtime="00:01:06.89" resultid="1306" heatid="2075" lane="4" entrytime="00:01:07.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="386" swimtime="00:01:15.92" resultid="1307" heatid="2104" lane="1" entrytime="00:01:15.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="420" swimtime="00:00:29.04" resultid="1308" heatid="2113" lane="5" />
                <RESULT eventid="1265" points="375" swimtime="00:00:27.95" resultid="1309" heatid="2133" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Poletti Veiga" birthdate="2010-10-01" gender="F" nation="BRA" license="376951" swrid="5603895" athleteid="1292" externalid="376951">
              <RESULTS>
                <RESULT eventid="1066" points="376" swimtime="00:02:48.78" resultid="1293" heatid="2042" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                    <SPLIT distance="100" swimtime="00:01:18.62" />
                    <SPLIT distance="150" swimtime="00:02:10.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1134" points="275" swimtime="00:01:23.02" resultid="1294" heatid="2073" lane="1" entrytime="00:01:19.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="497" swimtime="00:04:51.94" resultid="1295" heatid="2093" lane="3" entrytime="00:04:56.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                    <SPLIT distance="100" swimtime="00:01:10.99" />
                    <SPLIT distance="150" swimtime="00:01:48.11" />
                    <SPLIT distance="200" swimtime="00:02:25.62" />
                    <SPLIT distance="250" swimtime="00:03:02.66" />
                    <SPLIT distance="300" swimtime="00:03:39.99" />
                    <SPLIT distance="350" swimtime="00:04:17.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="345" swimtime="00:00:34.73" resultid="1296" heatid="2111" lane="3" entrytime="00:00:33.50" entrycourse="SCM" />
                <RESULT eventid="1260" points="465" swimtime="00:00:29.59" resultid="1297" heatid="2132" lane="4" entrytime="00:00:29.62" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco" lastname="Silva Telles" birthdate="2011-07-19" gender="M" nation="BRA" license="377311" swrid="5603911" athleteid="1310" externalid="377311">
              <RESULTS>
                <RESULT eventid="1070" points="211" swimtime="00:03:04.06" resultid="1311" heatid="2044" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.19" />
                    <SPLIT distance="100" swimtime="00:01:29.95" />
                    <SPLIT distance="150" swimtime="00:02:22.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="257" swimtime="00:00:39.24" resultid="1312" heatid="2085" lane="3" entrytime="00:00:43.37" entrycourse="SCM" />
                <RESULT eventid="1202" points="232" swimtime="00:01:29.87" resultid="1313" heatid="2103" lane="4" entrytime="00:01:37.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="243" swimtime="00:00:32.28" resultid="1314" heatid="2134" lane="3" entrytime="00:00:34.72" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Clara Bobroff" birthdate="2013-02-09" gender="F" nation="BRA" license="391752" swrid="5419807" athleteid="1315" externalid="391752">
              <RESULTS>
                <RESULT eventid="1077" points="225" swimtime="00:01:42.42" resultid="1316" heatid="2047" lane="5" entrytime="00:01:46.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="174" swimtime="00:00:45.19" resultid="1317" heatid="2056" lane="5" />
                <RESULT eventid="1144" points="300" swimtime="00:00:34.23" resultid="1318" heatid="2077" lane="4" entrytime="00:00:36.74" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Bordini Zocco" birthdate="2008-08-04" gender="F" nation="BRA" license="385677" swrid="5332871" athleteid="1282" externalid="385677">
              <RESULTS>
                <RESULT eventid="1083" points="359" swimtime="00:01:10.70" resultid="1283" heatid="2051" lane="5" entrytime="00:01:09.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1150" points="288" swimtime="00:00:42.92" resultid="1284" heatid="2082" lane="4" />
                <RESULT eventid="1134" points="304" swimtime="00:01:20.36" resultid="1285" heatid="2073" lane="6" entrytime="00:01:20.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="309" swimtime="00:01:32.18" resultid="1286" heatid="2102" lane="2" entrytime="00:01:30.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1241" points="295" swimtime="00:01:22.40" resultid="1287" heatid="2123" lane="2" entrytime="00:01:20.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Takemura Couto" birthdate="2010-02-08" gender="F" nation="BRA" license="376950" swrid="5603919" athleteid="1298" externalid="376950">
              <RESULTS>
                <RESULT eventid="1066" points="320" swimtime="00:02:58.04" resultid="1299" heatid="2042" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                    <SPLIT distance="100" swimtime="00:01:22.28" />
                    <SPLIT distance="150" swimtime="00:02:16.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1134" points="278" swimtime="00:01:22.75" resultid="1300" heatid="2073" lane="5" entrytime="00:01:18.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="373" swimtime="00:05:21.30" resultid="1301" heatid="2093" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                    <SPLIT distance="100" swimtime="00:01:13.87" />
                    <SPLIT distance="150" swimtime="00:01:54.12" />
                    <SPLIT distance="200" swimtime="00:02:34.72" />
                    <SPLIT distance="250" swimtime="00:03:15.56" />
                    <SPLIT distance="300" swimtime="00:03:57.28" />
                    <SPLIT distance="350" swimtime="00:04:39.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="422" swimtime="00:00:32.48" resultid="1302" heatid="2110" lane="2" />
                <RESULT eventid="1260" points="472" swimtime="00:00:29.45" resultid="1303" heatid="2132" lane="3" entrytime="00:00:29.14" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benjamin" lastname="Rinaldi Batistao" birthdate="2010-07-13" gender="M" nation="BRA" license="407035" swrid="5737920" athleteid="1325" externalid="407035">
              <RESULTS>
                <RESULT eventid="1091" points="271" swimtime="00:01:09.25" resultid="1326" heatid="2053" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="244" swimtime="00:00:34.76" resultid="1327" heatid="2113" lane="4" />
                <RESULT eventid="1265" points="274" swimtime="00:00:31.02" resultid="1328" heatid="2135" lane="6" entrytime="00:00:32.76" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Kikuchi Fujii" birthdate="2007-01-04" gender="M" nation="BRA" license="297805" swrid="5603863" athleteid="1276" externalid="297805" level="G-OLIMPICA">
              <RESULTS>
                <RESULT eventid="1070" points="610" swimtime="00:02:09.24" resultid="1277" heatid="2044" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.22" />
                    <SPLIT distance="100" swimtime="00:01:00.92" />
                    <SPLIT distance="150" swimtime="00:01:38.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1126" points="501" swimtime="00:00:27.83" resultid="1278" heatid="2067" lane="2" />
                <RESULT eventid="1157" points="570" swimtime="00:00:30.08" resultid="1279" heatid="2086" lane="4" entrytime="00:00:30.57" entrycourse="SCM" />
                <RESULT eventid="1202" points="666" swimtime="00:01:03.29" resultid="1280" heatid="2104" lane="3" entrytime="00:01:05.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="506" swimtime="00:01:00.65" resultid="1281" heatid="2125" lane="3" entrytime="00:01:01.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2864" nation="BRA" region="PR" clubid="1329" swrid="93756" name="Associacao De Pais E Amigos Da Natacao De Ponta Gr" shortname="Apan Ponta Grossa">
          <ATHLETES>
            <ATHLETE firstname="Sofia" lastname="Pontes Mattioli" birthdate="2011-09-10" gender="F" nation="BRA" license="366914" swrid="5602572" athleteid="1330" externalid="366914">
              <RESULTS>
                <RESULT eventid="1066" status="DNS" swimtime="00:00:00.00" resultid="1331" heatid="2042" lane="4" entrytime="00:03:03.97" entrycourse="SCM" />
                <RESULT eventid="1120" status="DNS" swimtime="00:00:00.00" resultid="1332" heatid="2066" lane="2" entrytime="00:00:37.97" entrycourse="SCM" />
                <RESULT eventid="1175" status="DNS" swimtime="00:00:00.00" resultid="1333" heatid="2093" lane="1" />
                <RESULT eventid="1219" status="DNS" swimtime="00:00:00.00" resultid="1334" heatid="2111" lane="5" entrytime="00:00:39.15" entrycourse="SCM" />
                <RESULT eventid="1241" status="DNS" swimtime="00:00:00.00" resultid="1335" heatid="2123" lane="6" entrytime="00:01:24.89" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18151" nation="BRA" region="PR" clubid="1600" swrid="95180" name="Clube Uniao Recreativo Palmense" shortname="Clube União">
          <ATHLETES>
            <ATHLETE firstname="Luiza" lastname="Langaro Spaniol" birthdate="2013-06-18" gender="F" nation="BRA" license="406600" swrid="5074027" athleteid="1601" externalid="406600">
              <RESULTS>
                <RESULT eventid="1077" points="344" swimtime="00:01:28.92" resultid="1602" heatid="2047" lane="4" entrytime="00:01:29.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="327" swimtime="00:00:36.64" resultid="1603" heatid="2057" lane="3" entrytime="00:00:37.45" entrycourse="SCM" />
                <RESULT eventid="1144" points="367" swimtime="00:00:32.00" resultid="1604" heatid="2078" lane="3" entrytime="00:00:32.09" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16053" nation="BRA" region="PR" clubid="1605" swrid="93777" name="Fábrica De Nadadores" shortname="Fábrica">
          <ATHLETES>
            <ATHLETE firstname="Dante" lastname="Gabriel Rossi" birthdate="2016-01-19" gender="M" nation="BRA" license="406928" swrid="5718627" athleteid="1775" externalid="406928">
              <RESULTS>
                <RESULT eventid="1167" points="71" swimtime="00:00:23.73" resultid="1776" heatid="2088" lane="3" entrytime="00:00:27.36" entrycourse="SCM" />
                <RESULT eventid="1188" points="71" swimtime="00:00:24.81" resultid="1777" heatid="2098" lane="5" />
                <RESULT eventid="1233" points="83" swimtime="00:00:46.06" resultid="1778" heatid="2116" lane="3" entrytime="00:00:58.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elen" lastname="Torres Gomes" birthdate="2015-10-15" gender="F" nation="BRA" license="396850" swrid="5641777" athleteid="1736" externalid="396850">
              <RESULTS>
                <RESULT eventid="1213" points="98" swimtime="00:00:54.72" resultid="1737" heatid="2108" lane="5" entrytime="00:00:52.93" entrycourse="SCM" />
                <RESULT eventid="1235" points="64" swimtime="00:01:10.58" resultid="1738" heatid="2118" lane="1" entrytime="00:01:10.06" entrycourse="SCM" />
                <RESULT eventid="1254" points="68" swimtime="00:00:56.07" resultid="1739" heatid="2127" lane="4" entrytime="00:00:52.88" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Bilemjian Leszczynski" birthdate="2014-02-22" gender="M" nation="BRA" license="406924" swrid="5631285" athleteid="1763" externalid="406924">
              <RESULTS>
                <RESULT eventid="1172" points="115" swimtime="00:01:32.13" resultid="1764" heatid="2091" lane="5" entrytime="00:01:51.25" entrycourse="SCM" />
                <RESULT eventid="1238" points="83" swimtime="00:00:57.18" resultid="1765" heatid="2120" lane="6" entrytime="00:00:59.86" entrycourse="SCM" />
                <RESULT eventid="1257" points="101" swimtime="00:00:43.27" resultid="1766" heatid="2130" lane="5" entrytime="00:00:48.21" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Dias Hei" birthdate="2016-01-22" gender="F" nation="BRA" license="414653" athleteid="1796" externalid="414653">
              <RESULTS>
                <RESULT eventid="1165" points="49" swimtime="00:00:30.38" resultid="1797" heatid="2087" lane="3" />
                <RESULT eventid="1186" points="49" swimtime="00:00:32.43" resultid="1798" heatid="2097" lane="1" />
                <RESULT eventid="1231" points="46" swimtime="00:01:03.87" resultid="1799" heatid="2115" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Kenji Yamaguchi" birthdate="2011-08-25" gender="M" nation="BRA" license="385708" swrid="5603862" athleteid="1666" externalid="385708">
              <RESULTS>
                <RESULT eventid="1070" points="247" swimtime="00:02:54.66" resultid="1667" heatid="2045" lane="6" entrytime="00:02:56.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                    <SPLIT distance="100" swimtime="00:01:20.75" />
                    <SPLIT distance="150" swimtime="00:02:12.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="181" swimtime="00:24:55.06" resultid="1668" heatid="2062" lane="3" />
                <RESULT eventid="1140" points="243" swimtime="00:01:16.51" resultid="1669" heatid="2075" lane="5" entrytime="00:01:14.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="165" swimtime="00:06:26.39" resultid="1670" heatid="2095" lane="4" />
                <RESULT eventid="1225" points="262" swimtime="00:00:33.98" resultid="1671" heatid="2114" lane="5" entrytime="00:00:34.85" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Souza" birthdate="2013-09-11" gender="M" nation="BRA" license="382211" swrid="5603916" athleteid="1752" externalid="382211">
              <RESULTS>
                <RESULT eventid="1063" points="184" swimtime="00:02:54.52" resultid="1753" heatid="2041" lane="2" entrytime="00:02:54.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.43" />
                    <SPLIT distance="100" swimtime="00:01:20.82" />
                    <SPLIT distance="150" swimtime="00:02:07.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="110" swimtime="00:01:39.54" resultid="1754" heatid="2065" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="183" swimtime="00:00:35.47" resultid="1755" heatid="2081" lane="1" entrytime="00:00:36.26" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Dias Rezende" birthdate="2016-03-04" gender="F" nation="BRA" license="406929" swrid="5631410" athleteid="1779" externalid="406929">
              <RESULTS>
                <RESULT eventid="1186" points="46" swimtime="00:00:32.97" resultid="1780" heatid="2097" lane="2" />
                <RESULT eventid="1209" points="30" swimtime="00:00:42.11" resultid="1781" heatid="2105" lane="4" />
                <RESULT eventid="1231" points="30" swimtime="00:01:13.22" resultid="1782" heatid="2115" lane="4" entrytime="00:01:24.31" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Livia" lastname="Eloisa Silva" birthdate="2012-03-03" gender="F" nation="BRA" license="399725" swrid="5651341" athleteid="1740" externalid="399725">
              <RESULTS>
                <RESULT eventid="1060" status="DNS" swimtime="00:00:00.00" resultid="1741" heatid="2038" lane="4" />
                <RESULT eventid="1099" status="DNS" swimtime="00:00:00.00" resultid="1742" heatid="2056" lane="2" entrytime="00:00:50.69" entrycourse="SCM" />
                <RESULT eventid="1144" status="DNS" swimtime="00:00:00.00" resultid="1743" heatid="2076" lane="5" entrytime="00:00:45.25" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Britto" birthdate="2012-10-04" gender="M" nation="BRA" license="378350" swrid="5588566" athleteid="1632" externalid="378350">
              <RESULTS>
                <RESULT eventid="1063" points="260" swimtime="00:02:35.57" resultid="1633" heatid="2041" lane="5" entrytime="00:02:54.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                    <SPLIT distance="100" swimtime="00:01:14.48" />
                    <SPLIT distance="150" swimtime="00:01:56.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1080" points="162" swimtime="00:01:41.22" resultid="1634" heatid="2049" lane="2" entrytime="00:01:40.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="176" swimtime="00:01:25.20" resultid="1635" heatid="2065" lane="3" entrytime="00:01:37.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Stephany" birthdate="2012-07-27" gender="F" nation="BRA" license="382210" swrid="5603917" athleteid="1756" externalid="382210">
              <RESULTS>
                <RESULT eventid="1060" points="235" swimtime="00:02:58.54" resultid="1757" heatid="2038" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                    <SPLIT distance="100" swimtime="00:01:26.52" />
                    <SPLIT distance="150" swimtime="00:02:13.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="145" swimtime="00:01:42.70" resultid="1758" heatid="2063" lane="5" entrytime="00:01:57.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1128" points="171" swimtime="00:03:39.23" resultid="1759" heatid="2069" lane="5" entrytime="00:03:38.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.00" />
                    <SPLIT distance="100" swimtime="00:01:44.56" />
                    <SPLIT distance="150" swimtime="00:02:50.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Rezende" birthdate="2012-01-23" gender="F" nation="BRA" license="370669" swrid="5603899" athleteid="1698" externalid="370669">
              <RESULTS>
                <RESULT eventid="1060" points="284" swimtime="00:02:47.77" resultid="1699" heatid="2039" lane="3" entrytime="00:02:49.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                    <SPLIT distance="100" swimtime="00:01:18.84" />
                    <SPLIT distance="150" swimtime="00:02:03.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="170" swimtime="00:01:52.51" resultid="1700" heatid="2047" lane="1" entrytime="00:02:02.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="260" swimtime="00:00:35.89" resultid="1701" heatid="2078" lane="6" entrytime="00:00:35.23" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monique" lastname="Istake" birthdate="2012-04-03" gender="F" nation="BRA" license="372023" swrid="5603857" athleteid="1636" externalid="372023">
              <RESULTS>
                <RESULT eventid="1077" status="DNS" swimtime="00:00:00.00" resultid="1637" heatid="2046" lane="2" />
                <RESULT eventid="1128" status="DNS" swimtime="00:00:00.00" resultid="1638" heatid="2069" lane="4" entrytime="00:03:07.98" entrycourse="SCM" />
                <RESULT eventid="1144" status="DNS" swimtime="00:00:00.00" resultid="1639" heatid="2078" lane="2" entrytime="00:00:34.12" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alex" lastname="Junior" birthdate="2013-03-11" gender="M" nation="BRA" license="385710" swrid="5603860" athleteid="1714" externalid="385710">
              <RESULTS>
                <RESULT eventid="1063" points="73" swimtime="00:03:56.78" resultid="1715" heatid="2040" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.71" />
                    <SPLIT distance="100" swimtime="00:01:48.02" />
                    <SPLIT distance="150" swimtime="00:02:53.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="62" swimtime="00:00:55.64" resultid="1716" heatid="2058" lane="2" />
                <RESULT eventid="1147" points="100" swimtime="00:00:43.38" resultid="1717" heatid="2079" lane="2" entrytime="00:00:46.98" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Gevaerd Verssutti Garcia" birthdate="2013-10-15" gender="F" nation="BRA" license="378404" swrid="5588723" athleteid="1702" externalid="378404">
              <RESULTS>
                <RESULT eventid="1099" points="253" swimtime="00:00:39.90" resultid="1703" heatid="2057" lane="5" entrytime="00:00:42.32" entrycourse="SCM" />
                <RESULT eventid="1128" points="217" swimtime="00:03:22.58" resultid="1704" heatid="2069" lane="6" entrytime="00:03:41.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.11" />
                    <SPLIT distance="100" swimtime="00:01:36.45" />
                    <SPLIT distance="150" swimtime="00:02:38.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="241" swimtime="00:00:36.82" resultid="1705" heatid="2077" lane="5" entrytime="00:00:38.72" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Limonta Moreto" birthdate="2015-06-29" gender="M" nation="BRA" license="408979" athleteid="1794" externalid="408979">
              <RESULTS>
                <RESULT eventid="1257" status="DNS" swimtime="00:00:00.00" resultid="1795" heatid="2129" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Pazinato" birthdate="2011-01-05" gender="M" nation="BRA" license="368149" swrid="5603889" athleteid="1672" externalid="368149">
              <RESULTS>
                <RESULT eventid="1109" points="268" swimtime="00:21:52.29" resultid="1673" heatid="2062" lane="2" />
                <RESULT eventid="1091" points="304" swimtime="00:01:06.63" resultid="1674" heatid="2054" lane="3" entrytime="00:01:06.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="280" swimtime="00:05:24.13" resultid="1675" heatid="2096" lane="6" entrytime="00:05:30.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.78" />
                    <SPLIT distance="100" swimtime="00:01:15.84" />
                    <SPLIT distance="150" swimtime="00:01:57.17" />
                    <SPLIT distance="200" swimtime="00:02:38.63" />
                    <SPLIT distance="250" swimtime="00:03:20.16" />
                    <SPLIT distance="300" swimtime="00:04:02.13" />
                    <SPLIT distance="350" swimtime="00:04:44.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="219" swimtime="00:01:20.16" resultid="1676" heatid="2125" lane="6" entrytime="00:01:18.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="285" swimtime="00:00:30.60" resultid="1677" heatid="2135" lane="5" entrytime="00:00:29.74" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Jupi Takaki" birthdate="2013-03-26" gender="F" nation="BRA" license="391845" swrid="5603861" athleteid="1718" externalid="391845">
              <RESULTS>
                <RESULT eventid="1060" points="274" swimtime="00:02:49.76" resultid="1719" heatid="2039" lane="5" entrytime="00:03:04.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.11" />
                    <SPLIT distance="100" swimtime="00:01:21.08" />
                    <SPLIT distance="150" swimtime="00:02:05.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="213" swimtime="00:01:30.42" resultid="1720" heatid="2063" lane="4" entrytime="00:01:35.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1128" points="218" swimtime="00:03:22.47" resultid="1721" heatid="2068" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.09" />
                    <SPLIT distance="100" swimtime="00:01:36.15" />
                    <SPLIT distance="150" swimtime="00:02:36.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruna" lastname="Scalise Drapzichinski" birthdate="2012-03-07" gender="F" nation="BRA" license="378349" swrid="5603909" athleteid="1618" externalid="378349">
              <RESULTS>
                <RESULT eventid="1077" points="430" swimtime="00:01:22.58" resultid="1619" heatid="2047" lane="3" entrytime="00:01:25.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1128" status="DNS" swimtime="00:00:00.00" resultid="1620" heatid="2069" lane="3" entrytime="00:03:07.73" entrycourse="SCM" />
                <RESULT eventid="1144" points="422" swimtime="00:00:30.55" resultid="1621" heatid="2078" lane="4" entrytime="00:00:32.43" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andressa" lastname="Zamarian Gouvea" birthdate="2007-09-18" gender="F" nation="BRA" license="318503" swrid="5603929" athleteid="1606" externalid="318503">
              <RESULTS>
                <RESULT eventid="1120" points="389" swimtime="00:00:34.57" resultid="1607" heatid="2066" lane="4" entrytime="00:00:34.98" entrycourse="SCM" />
                <RESULT eventid="1105" points="363" swimtime="00:21:13.00" resultid="1608" heatid="2060" lane="2" entrytime="00:21:46.88" entrycourse="SCM" />
                <RESULT eventid="1175" points="392" swimtime="00:05:15.81" resultid="1609" heatid="2093" lane="2" entrytime="00:05:16.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                    <SPLIT distance="100" swimtime="00:01:14.09" />
                    <SPLIT distance="150" swimtime="00:01:54.22" />
                    <SPLIT distance="200" swimtime="00:02:35.18" />
                    <SPLIT distance="250" swimtime="00:03:15.53" />
                    <SPLIT distance="300" swimtime="00:03:56.18" />
                    <SPLIT distance="350" swimtime="00:04:37.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="359" swimtime="00:00:34.28" resultid="1610" heatid="2111" lane="4" entrytime="00:00:33.90" entrycourse="SCM" />
                <RESULT eventid="1241" points="338" swimtime="00:01:18.73" resultid="1611" heatid="2123" lane="4" entrytime="00:01:16.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Bilemjian Leszczynski" birthdate="2011-08-06" gender="M" nation="BRA" license="406925" swrid="5587326" athleteid="1767" externalid="406925">
              <RESULTS>
                <RESULT eventid="1180" points="157" swimtime="00:06:32.97" resultid="1768" heatid="2094" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.73" />
                    <SPLIT distance="100" swimtime="00:01:27.99" />
                    <SPLIT distance="150" swimtime="00:02:17.23" />
                    <SPLIT distance="200" swimtime="00:03:06.61" />
                    <SPLIT distance="250" swimtime="00:03:58.20" />
                    <SPLIT distance="300" swimtime="00:04:50.30" />
                    <SPLIT distance="350" swimtime="00:05:41.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="113" swimtime="00:00:44.90" resultid="1769" heatid="2113" lane="3" />
                <RESULT eventid="1265" points="178" swimtime="00:00:35.79" resultid="1770" heatid="2134" lane="2" entrytime="00:00:36.56" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Traci Rodrigues" birthdate="2011-03-06" gender="M" nation="BRA" license="406927" swrid="5718893" athleteid="1622" externalid="406927">
              <RESULTS>
                <RESULT eventid="1091" status="DNS" swimtime="00:00:00.00" resultid="1623" heatid="2052" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:16.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" status="DNS" swimtime="00:00:00.00" resultid="1624" heatid="2084" lane="4" />
                <RESULT eventid="1180" points="135" swimtime="00:06:52.88" resultid="1625" heatid="2094" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.41" />
                    <SPLIT distance="100" swimtime="00:01:30.65" />
                    <SPLIT distance="150" swimtime="00:02:22.62" />
                    <SPLIT distance="200" swimtime="00:03:17.10" />
                    <SPLIT distance="250" swimtime="00:04:12.86" />
                    <SPLIT distance="300" swimtime="00:05:07.81" />
                    <SPLIT distance="350" swimtime="00:06:02.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="171" swimtime="00:01:39.51" resultid="1626" heatid="2103" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="204" swimtime="00:00:34.20" resultid="1627" heatid="2134" lane="5" entrytime="00:00:37.34" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Dias Rezende" birthdate="2016-03-04" gender="F" nation="BRA" license="406930" swrid="5685657" athleteid="1783" externalid="406930">
              <RESULTS>
                <RESULT eventid="1186" points="40" swimtime="00:00:34.47" resultid="1784" heatid="2097" lane="3" />
                <RESULT eventid="1209" points="73" swimtime="00:00:31.51" resultid="1785" heatid="2105" lane="2" />
                <RESULT eventid="1231" points="30" swimtime="00:01:13.20" resultid="1786" heatid="2115" lane="3" entrytime="00:01:13.75" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Magalhães Rezende" birthdate="2010-05-29" gender="F" nation="BRA" license="366960" swrid="5588793" athleteid="1650" externalid="366960">
              <RESULTS>
                <RESULT eventid="1083" points="359" swimtime="00:01:10.70" resultid="1651" heatid="2050" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="290" swimtime="00:22:51.69" resultid="1652" heatid="2060" lane="3" entrytime="00:22:31.63" entrycourse="SCM" />
                <RESULT eventid="1175" points="322" swimtime="00:05:37.43" resultid="1653" heatid="2093" lane="5" entrytime="00:05:34.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.21" />
                    <SPLIT distance="100" swimtime="00:01:14.96" />
                    <SPLIT distance="150" swimtime="00:01:57.03" />
                    <SPLIT distance="200" swimtime="00:02:39.46" />
                    <SPLIT distance="250" swimtime="00:03:23.14" />
                    <SPLIT distance="300" swimtime="00:04:07.88" />
                    <SPLIT distance="350" swimtime="00:04:53.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1241" points="309" swimtime="00:01:21.15" resultid="1654" heatid="2122" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1260" points="323" swimtime="00:00:33.41" resultid="1655" heatid="2132" lane="5" entrytime="00:00:31.73" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eloah" lastname="Juvedi Trindade" birthdate="2011-03-05" gender="F" nation="BRA" license="396829" swrid="5641768" athleteid="1728" externalid="396829">
              <RESULTS>
                <RESULT eventid="1066" points="197" swimtime="00:03:29.21" resultid="1729" heatid="2042" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.73" />
                    <SPLIT distance="100" swimtime="00:01:38.16" />
                    <SPLIT distance="150" swimtime="00:02:39.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1134" points="129" swimtime="00:01:46.90" resultid="1730" heatid="2072" lane="2" entrytime="00:01:50.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="242" swimtime="00:24:16.94" resultid="1731" heatid="2060" lane="1" />
                <RESULT eventid="1175" points="231" swimtime="00:06:16.94" resultid="1732" heatid="2092" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.26" />
                    <SPLIT distance="100" swimtime="00:01:22.98" />
                    <SPLIT distance="150" swimtime="00:02:10.74" />
                    <SPLIT distance="200" swimtime="00:03:01.11" />
                    <SPLIT distance="250" swimtime="00:03:52.87" />
                    <SPLIT distance="300" swimtime="00:04:43.23" />
                    <SPLIT distance="350" swimtime="00:05:31.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1241" points="229" swimtime="00:01:29.60" resultid="1733" heatid="2122" lane="3" entrytime="00:01:30.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Kuhnen Consalter" birthdate="2014-04-25" gender="F" nation="BRA" license="415372" athleteid="1800" externalid="415372">
              <RESULTS>
                <RESULT eventid="1254" points="172" swimtime="00:00:41.17" resultid="1801" heatid="2126" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Azevedo Martins" birthdate="2014-07-05" gender="F" nation="BRA" license="401859" swrid="5661340" athleteid="1744" externalid="401859">
              <RESULTS>
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="1745" heatid="2099" lane="3" entrytime="00:01:06.12" entrycourse="SCM" />
                <RESULT eventid="1235" status="DNS" swimtime="00:00:00.00" resultid="1746" heatid="2118" lane="2" entrytime="00:01:03.64" entrycourse="SCM" />
                <RESULT eventid="1254" status="DNS" swimtime="00:00:00.00" resultid="1747" heatid="2127" lane="2" entrytime="00:00:56.14" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Traci Rodrigues" birthdate="2014-10-27" gender="M" nation="BRA" license="406926" swrid="5726001" athleteid="1771" externalid="406926">
              <RESULTS>
                <RESULT eventid="1193" points="35" swimtime="00:01:06.36" resultid="1772" heatid="2101" lane="1" />
                <RESULT eventid="1238" points="89" swimtime="00:00:55.69" resultid="1773" heatid="2120" lane="2" entrytime="00:00:57.84" entrycourse="SCM" />
                <RESULT eventid="1257" points="108" swimtime="00:00:42.21" resultid="1774" heatid="2129" lane="3" entrytime="00:00:50.03" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Taparo" birthdate="2012-04-20" gender="F" nation="BRA" license="407283" swrid="5688565" athleteid="1790" externalid="407283">
              <RESULTS>
                <RESULT eventid="1099" status="DSQ" swimtime="00:00:46.05" resultid="1791" heatid="2056" lane="4" entrytime="00:00:45.66" entrycourse="SCM" />
                <RESULT eventid="1114" status="DSQ" swimtime="00:01:51.11" resultid="1792" heatid="2063" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="226" swimtime="00:00:37.59" resultid="1793" heatid="2077" lane="1" entrytime="00:00:39.33" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benicio" lastname="Garcia" birthdate="2011-09-09" gender="M" nation="BRA" license="378347" swrid="5603842" athleteid="1612" externalid="378347">
              <RESULTS>
                <RESULT eventid="1109" points="275" swimtime="00:21:41.50" resultid="1613" heatid="2062" lane="4" />
                <RESULT eventid="1091" points="234" swimtime="00:01:12.69" resultid="1614" heatid="2054" lane="2" entrytime="00:01:10.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="221" swimtime="00:05:50.90" resultid="1615" heatid="2095" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                    <SPLIT distance="100" swimtime="00:01:13.59" />
                    <SPLIT distance="150" swimtime="00:02:03.85" />
                    <SPLIT distance="200" swimtime="00:02:50.35" />
                    <SPLIT distance="250" swimtime="00:03:36.75" />
                    <SPLIT distance="300" swimtime="00:04:23.07" />
                    <SPLIT distance="350" swimtime="00:05:07.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" status="DNS" swimtime="00:00:00.00" resultid="1616" heatid="2114" lane="6" entrytime="00:00:37.70" entrycourse="SCM" />
                <RESULT eventid="1248" status="DNS" swimtime="00:00:00.00" resultid="1617" heatid="2125" lane="5" entrytime="00:01:17.15" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Ognibeni Paupitz" birthdate="2014-08-08" gender="F" nation="BRA" license="406923" swrid="5718889" athleteid="1760" externalid="406923">
              <RESULTS>
                <RESULT eventid="1235" points="118" swimtime="00:00:57.77" resultid="1761" heatid="2118" lane="5" entrytime="00:01:04.07" entrycourse="SCM" />
                <RESULT eventid="1254" points="139" swimtime="00:00:44.20" resultid="1762" heatid="2128" lane="1" entrytime="00:00:47.38" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Fernandes Dantas" birthdate="2016-12-14" gender="M" nation="BRA" license="406932" swrid="5700463" athleteid="1787" externalid="406932">
              <RESULTS>
                <RESULT eventid="1188" status="DNS" swimtime="00:00:00.00" resultid="1788" heatid="2098" lane="4" />
                <RESULT eventid="1233" status="DNS" swimtime="00:00:00.00" resultid="1789" heatid="2116" lane="2" entrytime="00:01:12.80" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Schmeiske Ruivo" birthdate="2013-10-21" gender="F" nation="BRA" license="402006" swrid="5661354" athleteid="1748" externalid="402006">
              <RESULTS>
                <RESULT eventid="1077" points="277" swimtime="00:01:35.62" resultid="1749" heatid="2047" lane="2" entrytime="00:01:40.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="227" swimtime="00:00:41.38" resultid="1750" heatid="2057" lane="4" entrytime="00:00:40.65" entrycourse="SCM" />
                <RESULT eventid="1144" points="315" swimtime="00:00:33.69" resultid="1751" heatid="2078" lane="5" entrytime="00:00:34.88" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Rossi" birthdate="2012-05-21" gender="M" nation="BRA" license="378346" swrid="5603901" athleteid="1690" externalid="378346">
              <RESULTS>
                <RESULT eventid="1063" points="236" swimtime="00:02:40.73" resultid="1691" heatid="2041" lane="4" entrytime="00:02:50.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                    <SPLIT distance="100" swimtime="00:01:16.38" />
                    <SPLIT distance="150" swimtime="00:01:58.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1080" points="142" swimtime="00:01:45.73" resultid="1692" heatid="2049" lane="5" entrytime="00:01:45.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="142" swimtime="00:01:31.53" resultid="1693" heatid="2065" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Lima Coelho" birthdate="2012-12-12" gender="M" nation="BRA" license="393775" swrid="5615959" athleteid="1640" externalid="393775">
              <RESULTS>
                <RESULT eventid="1063" points="141" swimtime="00:03:10.91" resultid="1641" heatid="2040" lane="3" entrytime="00:03:22.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.46" />
                    <SPLIT distance="100" swimtime="00:01:27.61" />
                    <SPLIT distance="150" swimtime="00:02:19.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="141" swimtime="00:00:42.43" resultid="1642" heatid="2059" lane="3" entrytime="00:00:42.35" entrycourse="SCM" />
                <RESULT eventid="1147" points="171" swimtime="00:00:36.31" resultid="1643" heatid="2080" lane="2" entrytime="00:00:38.30" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Silveira De Almeida" birthdate="2008-07-08" gender="M" nation="BRA" license="368152" swrid="5603912" athleteid="1678" externalid="368152">
              <RESULTS>
                <RESULT eventid="1070" points="361" swimtime="00:02:33.87" resultid="1679" heatid="2045" lane="4" entrytime="00:02:26.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.56" />
                    <SPLIT distance="100" swimtime="00:01:10.30" />
                    <SPLIT distance="150" swimtime="00:01:55.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="317" swimtime="00:01:10.05" resultid="1681" heatid="2075" lane="3" entrytime="00:01:01.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="272" swimtime="00:05:27.34" resultid="1682" heatid="2096" lane="4" entrytime="00:04:59.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.71" />
                    <SPLIT distance="100" swimtime="00:01:16.48" />
                    <SPLIT distance="150" swimtime="00:01:58.40" />
                    <SPLIT distance="200" swimtime="00:02:42.12" />
                    <SPLIT distance="250" swimtime="00:03:22.33" />
                    <SPLIT distance="300" swimtime="00:04:04.13" />
                    <SPLIT distance="350" swimtime="00:04:45.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" status="DNS" swimtime="00:00:00.00" resultid="1683" heatid="2124" lane="2" />
                <RESULT eventid="1109" points="242" swimtime="00:22:37.57" resultid="2145" heatid="2061" lane="5" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabel" lastname="Rezende" birthdate="2013-12-13" gender="F" nation="BRA" license="370657" swrid="5603900" athleteid="1628" externalid="370657">
              <RESULTS>
                <RESULT eventid="1077" points="143" swimtime="00:01:59.10" resultid="1629" heatid="2047" lane="6" entrytime="00:02:13.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1128" points="174" swimtime="00:03:38.27" resultid="1630" heatid="2068" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.74" />
                    <SPLIT distance="100" swimtime="00:01:46.19" />
                    <SPLIT distance="150" swimtime="00:02:51.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="230" swimtime="00:00:37.40" resultid="1631" heatid="2076" lane="2" entrytime="00:00:42.68" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Tiemi Yamaguchi" birthdate="2013-02-28" gender="F" nation="BRA" license="385707" swrid="5603920" athleteid="1706" externalid="385707">
              <RESULTS>
                <RESULT eventid="1099" points="222" swimtime="00:00:41.67" resultid="1707" heatid="2056" lane="6" />
                <RESULT eventid="1114" points="257" swimtime="00:01:25.00" resultid="1708" heatid="2063" lane="3" entrytime="00:01:26.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="276" swimtime="00:00:35.18" resultid="1709" heatid="2077" lane="6" entrytime="00:00:39.40" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Moreschi" birthdate="2012-08-09" gender="M" nation="BRA" license="385715" swrid="5603876" athleteid="1656" externalid="385715">
              <RESULTS>
                <RESULT eventid="1080" points="191" swimtime="00:01:35.84" resultid="1657" heatid="2049" lane="3" entrytime="00:01:34.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="140" swimtime="00:01:31.82" resultid="1658" heatid="2065" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="222" swimtime="00:00:33.29" resultid="1659" heatid="2081" lane="5" entrytime="00:00:35.48" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Bagatim" birthdate="2014-05-27" gender="F" nation="BRA" license="378353" swrid="5236649" athleteid="1694" externalid="378353">
              <RESULTS>
                <RESULT eventid="1169" points="235" swimtime="00:01:21.35" resultid="1695" heatid="2089" lane="3" entrytime="00:01:23.66" entrycourse="SCM" />
                <RESULT eventid="1190" points="240" swimtime="00:00:39.20" resultid="1696" heatid="2100" lane="3" entrytime="00:00:38.34" entrycourse="SCM" />
                <RESULT eventid="1213" points="173" swimtime="00:00:45.28" resultid="1697" heatid="2108" lane="2" entrytime="00:00:49.61" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theodoro" lastname="Marques Serra" birthdate="2009-11-24" gender="M" nation="BRA" license="370661" swrid="5603870" athleteid="1644" externalid="370661">
              <RESULTS>
                <RESULT eventid="1140" points="297" swimtime="00:01:11.59" resultid="1646" heatid="2074" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="404" swimtime="00:04:47.07" resultid="1647" heatid="2096" lane="2" entrytime="00:05:01.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                    <SPLIT distance="100" swimtime="00:01:06.60" />
                    <SPLIT distance="150" swimtime="00:01:43.84" />
                    <SPLIT distance="200" swimtime="00:02:21.06" />
                    <SPLIT distance="250" swimtime="00:02:58.47" />
                    <SPLIT distance="300" swimtime="00:03:35.28" />
                    <SPLIT distance="350" swimtime="00:04:11.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="372" swimtime="00:00:30.22" resultid="1648" heatid="2112" lane="2" />
                <RESULT eventid="1265" points="381" swimtime="00:00:27.79" resultid="1649" heatid="2135" lane="4" entrytime="00:00:29.22" entrycourse="SCM" />
                <RESULT eventid="1109" points="367" swimtime="00:19:42.61" resultid="2146" heatid="2061" lane="6" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Drapzichinski" birthdate="2015-08-21" gender="M" nation="BRA" license="391848" swrid="5603890" athleteid="1722" externalid="391848">
              <RESULTS>
                <RESULT eventid="1216" points="111" swimtime="00:00:45.94" resultid="1723" heatid="2109" lane="2" entrytime="00:00:51.97" entrycourse="SCM" />
                <RESULT eventid="1238" points="84" swimtime="00:00:56.86" resultid="1724" heatid="2119" lane="5" entrytime="00:01:09.38" entrycourse="SCM" />
                <RESULT eventid="1257" points="152" swimtime="00:00:37.75" resultid="1725" heatid="2130" lane="2" entrytime="00:00:42.94" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Valentina Gozaga" birthdate="2014-06-28" gender="F" nation="BRA" license="385709" swrid="5603924" athleteid="1710" externalid="385709">
              <RESULTS>
                <RESULT eventid="1169" status="DNS" swimtime="00:00:00.00" resultid="1711" heatid="2089" lane="4" entrytime="00:01:32.89" entrycourse="SCM" />
                <RESULT eventid="1213" status="DNS" swimtime="00:00:00.00" resultid="1712" heatid="2108" lane="4" entrytime="00:00:47.42" entrycourse="SCM" />
                <RESULT eventid="1254" status="DNS" swimtime="00:00:00.00" resultid="1713" heatid="2128" lane="3" entrytime="00:00:39.26" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="Jacobsen Donati" birthdate="2011-07-14" gender="M" nation="BRA" license="391851" swrid="5615735" athleteid="1660" externalid="391851">
              <RESULTS>
                <RESULT eventid="1070" status="DNS" swimtime="00:00:00.00" resultid="1661" heatid="2044" lane="3" entrytime="00:03:05.14" entrycourse="SCM" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="1662" heatid="2062" lane="5" />
                <RESULT eventid="1140" status="DNS" swimtime="00:00:00.00" resultid="1663" heatid="2075" lane="1" />
                <RESULT eventid="1180" status="DNS" swimtime="00:00:00.00" resultid="1664" heatid="2095" lane="3" entrytime="00:05:34.68" entrycourse="SCM" />
                <RESULT eventid="1265" points="345" swimtime="00:00:28.74" resultid="1665" heatid="2136" lane="1" entrytime="00:00:28.34" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Guinoza" birthdate="2013-01-06" gender="F" nation="BRA" license="392012" swrid="5510698" athleteid="1726" externalid="392012">
              <RESULTS>
                <RESULT eventid="1144" points="220" swimtime="00:00:37.98" resultid="1727" heatid="2076" lane="3" entrytime="00:00:39.92" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marco" lastname="Manzotti Marchi" birthdate="2015-06-26" gender="M" nation="BRA" license="396849" swrid="5641769" athleteid="1734" externalid="396849">
              <RESULTS>
                <RESULT eventid="1193" points="69" swimtime="00:00:52.83" resultid="1735" heatid="2101" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Braga" birthdate="2010-05-07" gender="M" nation="BRA" license="378345" swrid="5343953" athleteid="1684" externalid="378345">
              <RESULTS>
                <RESULT eventid="1070" points="347" swimtime="00:02:35.93" resultid="1685" heatid="2045" lane="5" entrytime="00:02:37.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.22" />
                    <SPLIT distance="100" swimtime="00:01:17.74" />
                    <SPLIT distance="150" swimtime="00:01:58.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="409" swimtime="00:00:33.59" resultid="1687" heatid="2086" lane="5" entrytime="00:00:33.67" entrycourse="SCM" />
                <RESULT eventid="1180" points="327" swimtime="00:05:07.82" resultid="1688" heatid="2096" lane="1" entrytime="00:05:07.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                    <SPLIT distance="100" swimtime="00:01:11.99" />
                    <SPLIT distance="150" swimtime="00:01:51.82" />
                    <SPLIT distance="200" swimtime="00:02:31.67" />
                    <SPLIT distance="250" swimtime="00:03:10.86" />
                    <SPLIT distance="300" swimtime="00:03:50.22" />
                    <SPLIT distance="350" swimtime="00:04:29.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="443" swimtime="00:01:12.47" resultid="1689" heatid="2104" lane="4" entrytime="00:01:13.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="297" swimtime="00:21:07.95" resultid="2144" heatid="2061" lane="4" late="yes" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2416" nation="BRA" region="PR" clubid="1336" swrid="93758" name="Apan/Maringá">
          <ATHLETES>
            <ATHLETE firstname="Pedro" lastname="Otavio Luz" birthdate="2013-07-27" gender="M" nation="BRA" license="392111" swrid="5603882" athleteid="1492" externalid="392111">
              <RESULTS>
                <RESULT eventid="1080" points="109" swimtime="00:01:55.71" resultid="1493" heatid="2048" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="169" swimtime="00:03:18.20" resultid="1494" heatid="2071" lane="3" entrytime="00:03:27.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.51" />
                    <SPLIT distance="100" swimtime="00:01:36.22" />
                    <SPLIT distance="150" swimtime="00:02:36.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="181" swimtime="00:00:35.59" resultid="1495" heatid="2080" lane="4" entrytime="00:00:36.95" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Antonio Mendes" birthdate="2008-12-04" gender="M" nation="BRA" license="366962" swrid="5196287" athleteid="1377" externalid="366962">
              <RESULTS>
                <RESULT eventid="1091" points="460" swimtime="00:00:58.08" resultid="1378" heatid="2052" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="505" swimtime="00:00:31.32" resultid="1379" heatid="2086" lane="2" entrytime="00:00:31.40" entrycourse="SCM" />
                <RESULT eventid="1265" status="DSQ" swimtime="00:00:25.61" resultid="1380" heatid="2136" lane="2" entrytime="00:00:26.95" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Bassil" birthdate="2015-07-02" gender="M" nation="BRA" license="407178" swrid="5718890" athleteid="1561" externalid="407178">
              <RESULTS>
                <RESULT eventid="1216" points="95" swimtime="00:00:48.44" resultid="1562" heatid="2109" lane="1" />
                <RESULT eventid="1238" points="85" swimtime="00:00:56.57" resultid="1563" heatid="2120" lane="1" entrytime="00:00:59.32" entrycourse="SCM" />
                <RESULT eventid="1257" points="101" swimtime="00:00:43.25" resultid="1564" heatid="2130" lane="1" entrytime="00:00:49.14" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raphael" lastname="Piai Pellegrini" birthdate="2012-03-24" gender="M" nation="BRA" license="377261" swrid="5603894" athleteid="1423" externalid="377261">
              <RESULTS>
                <RESULT eventid="1063" points="275" swimtime="00:02:32.77" resultid="1424" heatid="2041" lane="3" entrytime="00:02:24.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                    <SPLIT distance="100" swimtime="00:01:13.84" />
                    <SPLIT distance="150" swimtime="00:01:56.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="196" swimtime="00:03:08.42" resultid="1425" heatid="2070" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.96" />
                    <SPLIT distance="100" swimtime="00:01:24.99" />
                    <SPLIT distance="150" swimtime="00:02:26.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="250" swimtime="00:01:15.82" resultid="1426" heatid="2064" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Sanches Ghelere" birthdate="2008-08-06" gender="F" nation="BRA" license="372024" swrid="5603905" athleteid="1372" externalid="372024">
              <RESULTS>
                <RESULT eventid="1083" points="473" swimtime="00:01:04.46" resultid="1373" heatid="2051" lane="4" entrytime="00:01:04.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="392" swimtime="00:00:34.48" resultid="1374" heatid="2066" lane="3" entrytime="00:00:33.37" entrycourse="SCM" />
                <RESULT eventid="1175" points="438" swimtime="00:05:04.48" resultid="1375" heatid="2092" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.13" />
                    <SPLIT distance="100" swimtime="00:01:13.98" />
                    <SPLIT distance="150" swimtime="00:01:53.23" />
                    <SPLIT distance="200" swimtime="00:02:33.09" />
                    <SPLIT distance="250" swimtime="00:03:11.24" />
                    <SPLIT distance="300" swimtime="00:03:49.62" />
                    <SPLIT distance="350" swimtime="00:04:29.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="451" swimtime="00:00:31.78" resultid="1376" heatid="2110" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Eduardo Ebiner" birthdate="2013-07-29" gender="M" nation="BRA" license="397371" swrid="5641763" athleteid="1523" externalid="397371">
              <RESULTS>
                <RESULT eventid="1063" points="161" swimtime="00:03:02.46" resultid="1524" heatid="2040" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.52" />
                    <SPLIT distance="100" swimtime="00:01:27.84" />
                    <SPLIT distance="150" swimtime="00:02:15.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="96" swimtime="00:00:48.18" resultid="1525" heatid="2058" lane="4" />
                <RESULT eventid="1131" points="132" swimtime="00:03:35.25" resultid="1526" heatid="2070" lane="3" entrytime="00:03:50.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.78" />
                    <SPLIT distance="100" swimtime="00:01:48.57" />
                    <SPLIT distance="150" swimtime="00:02:48.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Peroni Passafaro" birthdate="2013-09-17" gender="F" nation="BRA" license="370659" swrid="5603893" athleteid="1400" externalid="370659">
              <RESULTS>
                <RESULT eventid="1077" points="154" swimtime="00:01:56.17" resultid="1401" heatid="2046" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="158" swimtime="00:01:39.96" resultid="1402" heatid="2063" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="240" swimtime="00:00:36.87" resultid="1403" heatid="2078" lane="1" entrytime="00:00:35.21" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Biason Santana" birthdate="2009-01-21" gender="M" nation="BRA" license="366969" swrid="5317765" athleteid="1381" externalid="366969">
              <RESULTS>
                <RESULT eventid="1091" points="443" swimtime="00:00:58.82" resultid="1382" heatid="2055" lane="4" entrytime="00:01:00.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="496" swimtime="00:00:27.47" resultid="1383" heatid="2114" lane="4" entrytime="00:00:28.15" entrycourse="SCM" />
                <RESULT eventid="1248" points="293" swimtime="00:01:12.74" resultid="1384" heatid="2124" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lara" lastname="Constantino" birthdate="2012-06-02" gender="F" nation="BRA" license="382208" swrid="5420069" athleteid="1439" externalid="382208">
              <RESULTS>
                <RESULT eventid="1060" points="210" swimtime="00:03:05.36" resultid="1440" heatid="2039" lane="2" entrytime="00:03:02.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.54" />
                    <SPLIT distance="100" swimtime="00:01:30.14" />
                    <SPLIT distance="150" swimtime="00:02:18.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="231" swimtime="00:00:41.10" resultid="1441" heatid="2056" lane="3" entrytime="00:00:45.37" entrycourse="SCM" />
                <RESULT eventid="1128" points="243" swimtime="00:03:15.07" resultid="1442" heatid="2069" lane="2" entrytime="00:03:36.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.86" />
                    <SPLIT distance="150" swimtime="00:02:28.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laion" lastname="Miguel Simoes" birthdate="2016-04-02" gender="M" nation="BRA" license="407179" swrid="5718695" athleteid="1565" externalid="407179">
              <RESULTS>
                <RESULT eventid="1167" points="50" swimtime="00:00:26.79" resultid="1566" heatid="2088" lane="4" entrytime="00:00:36.50" entrycourse="SCM" />
                <RESULT eventid="1188" points="49" swimtime="00:00:28.08" resultid="1567" heatid="2098" lane="3" entrytime="00:00:33.37" entrycourse="SCM" />
                <RESULT eventid="1211" points="66" swimtime="00:00:28.31" resultid="1568" heatid="2106" lane="3" entrytime="00:00:37.92" entrycourse="SCM" />
                <RESULT eventid="1233" points="55" swimtime="00:00:52.93" resultid="1569" heatid="2116" lane="4" entrytime="00:01:05.23" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Pacheco" birthdate="2012-10-03" gender="M" nation="BRA" license="370663" swrid="5603883" athleteid="1408" externalid="370663">
              <RESULTS>
                <RESULT eventid="1080" points="206" swimtime="00:01:33.45" resultid="1409" heatid="2048" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="188" swimtime="00:01:23.31" resultid="1410" heatid="2064" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="250" swimtime="00:00:31.97" resultid="1411" heatid="2081" lane="4" entrytime="00:00:31.96" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="De Desvars" birthdate="2016-04-08" gender="F" nation="BRA" license="414853" athleteid="1596" externalid="414853">
              <RESULTS>
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="1597" heatid="2087" lane="4" />
                <RESULT eventid="1186" status="DNS" swimtime="00:00:00.00" resultid="1598" heatid="2097" lane="5" />
                <RESULT eventid="1231" status="DNS" swimtime="00:00:00.00" resultid="1599" heatid="2115" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Allyce" lastname="Rodrigues Tavares" birthdate="2014-10-13" gender="F" nation="BRA" license="403389" swrid="5676291" athleteid="1543" externalid="403389">
              <RESULTS>
                <RESULT eventid="1213" points="31" swimtime="00:01:19.82" resultid="1544" heatid="2107" lane="4" entrytime="00:01:17.76" entrycourse="SCM" />
                <RESULT eventid="1254" points="20" swimtime="00:01:23.58" resultid="1545" heatid="2126" lane="3" entrytime="00:01:27.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Martins Pedro" birthdate="2015-01-19" gender="F" nation="BRA" license="403390" swrid="5676290" athleteid="1546" externalid="403390">
              <RESULTS>
                <RESULT eventid="1190" points="49" swimtime="00:01:06.45" resultid="1547" heatid="2100" lane="2" entrytime="00:01:02.78" entrycourse="SCM" />
                <RESULT eventid="1213" points="69" swimtime="00:01:01.46" resultid="1548" heatid="2107" lane="2" />
                <RESULT eventid="1254" points="91" swimtime="00:00:50.81" resultid="1549" heatid="2128" lane="6" entrytime="00:00:50.54" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Chaim" birthdate="2011-05-29" gender="F" nation="BRA" license="370662" swrid="5409721" athleteid="1404" externalid="370662">
              <RESULTS>
                <RESULT eventid="1083" points="309" swimtime="00:01:14.31" resultid="1405" heatid="2050" lane="3" entrytime="00:01:15.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="289" swimtime="00:05:49.65" resultid="1406" heatid="2092" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.51" />
                    <SPLIT distance="100" swimtime="00:01:20.06" />
                    <SPLIT distance="150" swimtime="00:02:04.00" />
                    <SPLIT distance="200" swimtime="00:02:49.83" />
                    <SPLIT distance="250" swimtime="00:03:35.09" />
                    <SPLIT distance="300" swimtime="00:04:20.40" />
                    <SPLIT distance="350" swimtime="00:05:05.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1241" points="243" swimtime="00:01:27.86" resultid="1407" heatid="2122" lane="4" entrytime="00:01:31.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Campos" birthdate="2013-02-17" gender="M" nation="BRA" license="377262" swrid="5641756" athleteid="1427" externalid="377262">
              <RESULTS>
                <RESULT eventid="1080" points="122" swimtime="00:01:51.28" resultid="1428" heatid="2048" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="93" swimtime="00:01:45.16" resultid="1429" heatid="2065" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="162" swimtime="00:00:36.95" resultid="1430" heatid="2081" lane="6" entrytime="00:00:36.40" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Otavio Costa" birthdate="2009-01-28" gender="M" nation="BRA" license="370666" swrid="5603881" athleteid="1412" externalid="370666">
              <RESULTS>
                <RESULT eventid="1140" points="218" swimtime="00:01:19.33" resultid="1413" heatid="2074" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="250" swimtime="00:00:39.58" resultid="1414" heatid="2084" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Rampasi" birthdate="2013-10-16" gender="F" nation="BRA" license="382209" swrid="5603866" athleteid="1443" externalid="382209">
              <RESULTS>
                <RESULT eventid="1060" points="198" swimtime="00:03:09.06" resultid="1444" heatid="2039" lane="1" entrytime="00:03:11.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.64" />
                    <SPLIT distance="100" swimtime="00:01:32.69" />
                    <SPLIT distance="150" swimtime="00:02:21.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="105" swimtime="00:00:53.42" resultid="1445" heatid="2056" lane="1" />
                <RESULT eventid="1128" points="178" swimtime="00:03:36.58" resultid="1446" heatid="2068" lane="3" entrytime="00:04:11.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.69" />
                    <SPLIT distance="100" swimtime="00:01:49.30" />
                    <SPLIT distance="150" swimtime="00:02:51.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Pastre" birthdate="2014-03-10" gender="F" nation="BRA" license="403760" swrid="5684593" athleteid="1550" externalid="403760">
              <RESULTS>
                <RESULT eventid="1190" points="142" swimtime="00:00:46.66" resultid="1551" heatid="2100" lane="5" entrytime="00:01:05.07" entrycourse="SCM" />
                <RESULT eventid="1213" points="244" swimtime="00:00:40.36" resultid="1552" heatid="2108" lane="3" entrytime="00:00:40.48" entrycourse="SCM" />
                <RESULT eventid="1254" points="204" swimtime="00:00:38.93" resultid="1553" heatid="2128" lane="4" entrytime="00:00:40.61" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Felipe Sakaguti" birthdate="2007-06-22" gender="M" nation="BRA" license="407187" swrid="5688778" athleteid="1578" externalid="407187">
              <RESULTS>
                <RESULT eventid="1091" status="DNS" swimtime="00:00:00.00" resultid="1579" heatid="2054" lane="6" entrytime="00:01:38.45" entrycourse="SCM" />
                <RESULT eventid="1126" status="DNS" swimtime="00:00:00.00" resultid="1580" heatid="2067" lane="4" entrytime="00:00:55.25" entrycourse="SCM" />
                <RESULT eventid="1265" points="105" swimtime="00:00:42.66" resultid="1581" heatid="2134" lane="1" entrytime="00:00:44.33" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Andrade Silva" birthdate="2016-03-15" gender="M" nation="BRA" license="414852" athleteid="1591" externalid="414852">
              <RESULTS>
                <RESULT eventid="1167" points="36" swimtime="00:00:29.82" resultid="1592" heatid="2088" lane="2" />
                <RESULT eventid="1188" points="90" swimtime="00:00:22.94" resultid="1593" heatid="2098" lane="2" />
                <RESULT eventid="1211" points="61" swimtime="00:00:29.11" resultid="1594" heatid="2106" lane="4" />
                <RESULT eventid="1233" points="79" swimtime="00:00:46.90" resultid="1595" heatid="2116" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Sol Reolon Gomes" birthdate="2011-02-28" gender="F" nation="BRA" license="392100" swrid="5603914" athleteid="1465" externalid="392100">
              <RESULTS>
                <RESULT eventid="1083" points="411" swimtime="00:01:07.57" resultid="1466" heatid="2051" lane="2" entrytime="00:01:08.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1241" points="376" swimtime="00:01:16.02" resultid="1467" heatid="2123" lane="5" entrytime="00:01:20.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Siqueira Almeida" birthdate="2016-06-21" gender="F" nation="BRA" license="414848" athleteid="1582" externalid="414848">
              <RESULTS>
                <RESULT eventid="1165" points="70" swimtime="00:00:27.07" resultid="1583" heatid="2087" lane="2" />
                <RESULT eventid="1186" points="92" swimtime="00:00:26.25" resultid="1584" heatid="2097" lane="4" />
                <RESULT eventid="1209" points="73" swimtime="00:00:31.49" resultid="1585" heatid="2105" lane="3" />
                <RESULT eventid="1231" points="59" swimtime="00:00:58.80" resultid="1586" heatid="2115" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wellington" lastname="De Lima" birthdate="2008-03-01" gender="M" nation="BRA" license="370024" swrid="5470912" athleteid="1344" externalid="370024">
              <RESULTS>
                <RESULT eventid="1265" points="461" swimtime="00:00:26.09" resultid="1345" heatid="2136" lane="4" entrytime="00:00:25.99" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heitor" lastname="Bello Paula" birthdate="2015-06-14" gender="M" nation="BRA" license="393776" swrid="5507529" athleteid="1511" externalid="393776">
              <RESULTS>
                <RESULT eventid="1172" points="98" swimtime="00:01:37.06" resultid="1512" heatid="2090" lane="2" />
                <RESULT eventid="1216" points="106" swimtime="00:00:46.58" resultid="1513" heatid="2109" lane="5" entrytime="00:00:56.00" entrycourse="SCM" />
                <RESULT eventid="1238" points="70" swimtime="00:01:00.40" resultid="1514" heatid="2119" lane="4" entrytime="00:01:02.70" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Muniz" birthdate="2012-09-03" gender="M" nation="BRA" license="392106" swrid="5603877" athleteid="1480" externalid="392106">
              <RESULTS>
                <RESULT eventid="1063" points="151" swimtime="00:03:06.52" resultid="1481" heatid="2040" lane="4" entrytime="00:03:37.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.72" />
                    <SPLIT distance="100" swimtime="00:01:33.50" />
                    <SPLIT distance="150" swimtime="00:02:23.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="98" swimtime="00:00:47.95" resultid="1482" heatid="2059" lane="4" entrytime="00:00:47.51" entrycourse="SCM" />
                <RESULT eventid="1147" points="184" swimtime="00:00:35.40" resultid="1483" heatid="2080" lane="1" entrytime="00:00:40.27" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Garcia Cavalcante" birthdate="2011-11-21" gender="M" nation="BRA" license="378200" swrid="5603840" athleteid="1353" externalid="378200">
              <RESULTS>
                <RESULT eventid="1140" points="149" swimtime="00:01:29.96" resultid="1354" heatid="2074" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="278" swimtime="00:01:24.65" resultid="1355" heatid="2103" lane="3" entrytime="00:01:25.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Isabel Henriques" birthdate="2007-09-05" gender="F" nation="BRA" license="414491" athleteid="1360" externalid="414491">
              <RESULTS>
                <RESULT eventid="1083" points="172" swimtime="00:01:30.33" resultid="1361" heatid="2050" lane="2" entrytime="00:01:33.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="135" swimtime="00:00:49.17" resultid="1362" heatid="2066" lane="1" entrytime="00:00:50.11" entrycourse="SCM" />
                <RESULT eventid="1260" points="179" swimtime="00:00:40.64" resultid="1363" heatid="2131" lane="3" entrytime="00:00:41.40" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Santos Carraro" birthdate="2014-06-04" gender="M" nation="BRA" license="392097" swrid="5603908" athleteid="1458" externalid="392097">
              <RESULTS>
                <RESULT eventid="1172" points="163" swimtime="00:01:21.97" resultid="1459" heatid="2091" lane="4" entrytime="00:01:24.90" entrycourse="SCM" />
                <RESULT eventid="1193" points="126" swimtime="00:00:43.34" resultid="1460" heatid="2101" lane="3" entrytime="00:00:45.43" entrycourse="SCM" />
                <RESULT eventid="1238" points="99" swimtime="00:00:53.87" resultid="1461" heatid="2119" lane="3" entrytime="00:01:00.65" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Arthur Da Silva Ortiz" birthdate="2015-04-20" gender="M" nation="BRA" license="399733" swrid="5676285" athleteid="1527" externalid="399733">
              <RESULTS>
                <RESULT eventid="1172" points="140" swimtime="00:01:26.35" resultid="1528" heatid="2090" lane="3" />
                <RESULT eventid="1193" points="89" swimtime="00:00:48.66" resultid="1529" heatid="2101" lane="2" entrytime="00:00:50.56" entrycourse="SCM" />
                <RESULT eventid="1238" points="110" swimtime="00:00:52.04" resultid="1530" heatid="2120" lane="3" entrytime="00:00:53.59" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Junio Brambilla" birthdate="2002-04-08" gender="M" nation="BRA" license="392112" swrid="5603859" athleteid="1496" externalid="392112">
              <RESULTS>
                <RESULT eventid="1225" points="319" swimtime="00:00:31.80" resultid="1497" heatid="2112" lane="3" />
                <RESULT eventid="1265" points="256" swimtime="00:00:31.73" resultid="1498" heatid="2134" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Furuchi Martins" birthdate="2011-10-05" gender="F" nation="BRA" license="367001" swrid="5602616" athleteid="1499" externalid="367001">
              <RESULTS>
                <RESULT eventid="1150" points="322" swimtime="00:00:41.37" resultid="1500" heatid="2083" lane="2" entrytime="00:00:44.08" entrycourse="SCM" />
                <RESULT eventid="1196" points="317" swimtime="00:01:31.44" resultid="1501" heatid="2102" lane="1" entrytime="00:01:34.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1241" points="212" swimtime="00:01:32.01" resultid="1502" heatid="2121" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juan" lastname="Bernardo Padua" birthdate="2013-07-15" gender="M" nation="BRA" license="392108" swrid="5305422" athleteid="1484" externalid="392108">
              <RESULTS>
                <RESULT eventid="1063" points="185" swimtime="00:02:54.32" resultid="1485" heatid="2041" lane="6" entrytime="00:03:08.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.72" />
                    <SPLIT distance="100" swimtime="00:01:21.19" />
                    <SPLIT distance="150" swimtime="00:02:09.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="141" swimtime="00:00:42.43" resultid="1486" heatid="2059" lane="5" />
                <RESULT eventid="1131" points="190" swimtime="00:03:10.63" resultid="1487" heatid="2071" lane="4" entrytime="00:03:29.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.36" />
                    <SPLIT distance="100" swimtime="00:01:34.94" />
                    <SPLIT distance="150" swimtime="00:02:27.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Passafaro" birthdate="2009-02-01" gender="F" nation="BRA" license="370673" swrid="5603885" athleteid="1369" externalid="370673">
              <RESULTS>
                <RESULT eventid="1134" points="275" swimtime="00:01:23.07" resultid="1370" heatid="2072" lane="3" entrytime="00:01:24.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1219" points="399" swimtime="00:00:33.10" resultid="1371" heatid="2111" lane="2" entrytime="00:00:34.72" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Batista Sanchez" birthdate="2009-05-22" gender="M" nation="BRA" license="370668" swrid="5255779" athleteid="1346" externalid="370668">
              <RESULTS>
                <RESULT eventid="1070" points="374" swimtime="00:02:32.12" resultid="1347" heatid="2044" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                    <SPLIT distance="100" swimtime="00:01:14.90" />
                    <SPLIT distance="150" swimtime="00:01:56.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="452" swimtime="00:01:11.99" resultid="1348" heatid="2104" lane="5" entrytime="00:01:14.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Pavão" birthdate="2012-04-04" gender="F" nation="BRA" license="377259" swrid="5603888" athleteid="1415" externalid="377259">
              <RESULTS>
                <RESULT eventid="1077" points="217" swimtime="00:01:43.62" resultid="1416" heatid="2046" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="234" swimtime="00:00:40.95" resultid="1417" heatid="2057" lane="2" entrytime="00:00:41.32" entrycourse="SCM" />
                <RESULT eventid="1144" points="297" swimtime="00:00:34.35" resultid="1418" heatid="2077" lane="3" entrytime="00:00:35.79" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carina" lastname="Costa Profeta" birthdate="2008-03-20" gender="F" nation="BRA" license="366964" swrid="5591584" athleteid="1364" externalid="366964">
              <RESULTS>
                <RESULT eventid="1196" points="464" swimtime="00:01:20.52" resultid="1365" heatid="2102" lane="3" entrytime="00:01:17.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felype" lastname="Gongora Zago" birthdate="2011-09-14" gender="M" nation="BRA" license="392099" swrid="5603848" athleteid="1462" externalid="392099">
              <RESULTS>
                <RESULT eventid="1091" points="214" swimtime="00:01:14.86" resultid="1463" heatid="2054" lane="1" entrytime="00:01:16.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="193" swimtime="00:00:37.63" resultid="1464" heatid="2114" lane="1" entrytime="00:00:35.97" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Catarina" lastname="Wendt Jesus" birthdate="2013-07-09" gender="F" nation="BRA" license="393778" swrid="5641780" athleteid="1515" externalid="393778">
              <RESULTS>
                <RESULT eventid="1060" points="337" swimtime="00:02:38.46" resultid="1516" heatid="2039" lane="4" entrytime="00:02:58.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                    <SPLIT distance="100" swimtime="00:01:16.26" />
                    <SPLIT distance="150" swimtime="00:01:58.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="291" swimtime="00:00:38.08" resultid="1517" heatid="2057" lane="1" entrytime="00:00:43.48" entrycourse="SCM" />
                <RESULT eventid="1114" points="268" swimtime="00:01:23.75" resultid="1518" heatid="2063" lane="2" entrytime="00:01:38.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Schuch Pimpao" birthdate="2010-05-17" gender="M" nation="BRA" license="355586" swrid="5588908" athleteid="1385" externalid="355586">
              <RESULTS>
                <RESULT eventid="1070" points="336" swimtime="00:02:37.59" resultid="1386" heatid="2045" lane="2" entrytime="00:02:34.86" entrycourse="SCM" />
                <RESULT eventid="1202" points="328" swimtime="00:01:20.12" resultid="1387" heatid="2104" lane="6" entrytime="00:01:21.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="317" swimtime="00:01:10.87" resultid="1388" heatid="2125" lane="4" entrytime="00:01:08.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietro" lastname="Nabas De Assis" birthdate="2011-07-09" gender="M" nation="BRA" license="366968" swrid="5603878" athleteid="1392" externalid="366968">
              <RESULTS>
                <RESULT eventid="1070" points="263" swimtime="00:02:51.03" resultid="1393" heatid="2045" lane="1" entrytime="00:02:53.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.76" />
                    <SPLIT distance="100" swimtime="00:01:23.07" />
                    <SPLIT distance="150" swimtime="00:02:10.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="283" swimtime="00:00:37.96" resultid="1394" heatid="2086" lane="1" entrytime="00:00:34.95" entrycourse="SCM" />
                <RESULT eventid="1180" points="289" swimtime="00:05:20.68" resultid="1395" heatid="2095" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.51" />
                    <SPLIT distance="100" swimtime="00:01:14.23" />
                    <SPLIT distance="150" swimtime="00:01:56.21" />
                    <SPLIT distance="200" swimtime="00:02:38.01" />
                    <SPLIT distance="250" swimtime="00:03:19.50" />
                    <SPLIT distance="300" swimtime="00:04:01.39" />
                    <SPLIT distance="350" swimtime="00:04:41.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Ayres" birthdate="2012-05-05" gender="M" nation="BRA" license="378035" swrid="5208079" athleteid="1431" externalid="378035">
              <RESULTS>
                <RESULT eventid="1080" points="194" swimtime="00:01:35.34" resultid="1432" heatid="2049" lane="4" entrytime="00:01:35.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="261" swimtime="00:01:14.70" resultid="1433" heatid="2064" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="276" swimtime="00:00:30.93" resultid="1434" heatid="2081" lane="3" entrytime="00:00:31.05" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Mendes Costa" birthdate="2014-04-03" gender="F" nation="BRA" license="378341" swrid="5603873" athleteid="1557" externalid="378341">
              <RESULTS>
                <RESULT eventid="1190" points="88" swimtime="00:00:54.80" resultid="1558" heatid="2100" lane="4" entrytime="00:00:54.62" entrycourse="SCM" />
                <RESULT eventid="1235" points="113" swimtime="00:00:58.65" resultid="1559" heatid="2118" lane="4" entrytime="00:00:58.27" entrycourse="SCM" />
                <RESULT eventid="1254" status="DNS" swimtime="00:00:00.00" resultid="1560" heatid="2128" lane="5" entrytime="00:00:45.47" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Marques" birthdate="2015-10-15" gender="F" nation="BRA" license="399738" swrid="5651346" athleteid="1531" externalid="399738">
              <RESULTS>
                <RESULT eventid="1213" points="40" swimtime="00:01:13.36" resultid="1532" heatid="2107" lane="3" entrytime="00:01:15.08" entrycourse="SCM" />
                <RESULT eventid="1235" points="26" swimtime="00:01:35.58" resultid="1533" heatid="2117" lane="3" entrytime="00:01:41.83" entrycourse="SCM" />
                <RESULT eventid="1254" points="27" swimtime="00:01:15.75" resultid="1534" heatid="2127" lane="1" entrytime="00:01:16.99" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Campelo" birthdate="2011-09-12" gender="M" nation="BRA" license="366963" swrid="5588742" athleteid="1389" externalid="366963">
              <RESULTS>
                <RESULT eventid="1091" points="444" swimtime="00:00:58.76" resultid="1390" heatid="2055" lane="5" entrytime="00:01:02.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="335" swimtime="00:01:09.57" resultid="1391" heatid="2125" lane="2" entrytime="00:01:13.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabrielle" lastname="Borba" birthdate="2014-06-15" gender="F" nation="BRA" license="385705" swrid="5323267" athleteid="1447" externalid="385705">
              <RESULTS>
                <RESULT eventid="1213" points="103" swimtime="00:00:53.78" resultid="1448" heatid="2108" lane="1" entrytime="00:00:55.49" entrycourse="SCM" />
                <RESULT eventid="1235" points="143" swimtime="00:00:54.15" resultid="1449" heatid="2118" lane="3" entrytime="00:00:57.94" entrycourse="SCM" />
                <RESULT eventid="1254" points="153" swimtime="00:00:42.84" resultid="1450" heatid="2128" lane="2" entrytime="00:00:44.25" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Ghelere" birthdate="2011-04-03" gender="F" nation="BRA" license="368146" swrid="5603843" athleteid="1396" externalid="368146">
              <RESULTS>
                <RESULT eventid="1083" points="312" swimtime="00:01:14.02" resultid="1397" heatid="2051" lane="1" entrytime="00:01:10.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1134" status="DSQ" swimtime="00:01:25.59" resultid="1398" heatid="2072" lane="4" entrytime="00:01:28.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1241" status="DSQ" swimtime="00:01:22.48" resultid="1399" heatid="2123" lane="1" entrytime="00:01:21.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Donato De Morais" birthdate="2009-03-28" gender="F" nation="BRA" license="345588" swrid="5485198" athleteid="1366" externalid="345588">
              <RESULTS>
                <RESULT eventid="1083" points="379" swimtime="00:01:09.41" resultid="1367" heatid="2051" lane="6" entrytime="00:01:11.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1241" points="386" swimtime="00:01:15.37" resultid="1368" heatid="2123" lane="3" entrytime="00:01:16.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lavinia" lastname="Bossoni" birthdate="2013-11-03" gender="F" nation="BRA" license="377260" swrid="5343093" athleteid="1419" externalid="377260">
              <RESULTS>
                <RESULT eventid="1077" points="199" swimtime="00:01:46.65" resultid="1420" heatid="2046" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1128" points="176" swimtime="00:03:37.05" resultid="1421" heatid="2069" lane="1" entrytime="00:03:39.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.22" />
                    <SPLIT distance="100" swimtime="00:01:47.13" />
                    <SPLIT distance="150" swimtime="00:02:49.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="202" swimtime="00:00:39.07" resultid="1422" heatid="2076" lane="4" entrytime="00:00:40.91" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Pauloski Murante" birthdate="1997-06-06" gender="M" nation="BRA" license="367086" swrid="5603887" athleteid="1554" externalid="367086">
              <RESULTS>
                <RESULT eventid="1091" points="277" swimtime="00:01:08.72" resultid="1555" heatid="2054" lane="5" entrytime="00:01:10.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1265" points="285" swimtime="00:00:30.60" resultid="1556" heatid="2133" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathan" lastname="Novak Pinho" birthdate="2012-11-14" gender="M" nation="BRA" license="378199" swrid="5603879" athleteid="1435" externalid="378199">
              <RESULTS>
                <RESULT eventid="1080" points="95" swimtime="00:02:01.12" resultid="1436" heatid="2049" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" status="DSQ" swimtime="00:03:24.29" resultid="1437" heatid="2070" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.89" />
                    <SPLIT distance="100" swimtime="00:01:31.20" />
                    <SPLIT distance="150" swimtime="00:02:40.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="207" swimtime="00:00:34.04" resultid="1438" heatid="2080" lane="3" entrytime="00:00:36.88" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnes" lastname="Sophie Amadei" birthdate="2014-01-10" gender="F" nation="BRA" license="403388" swrid="5676293" athleteid="1539" externalid="403388">
              <RESULTS>
                <RESULT eventid="1190" points="98" swimtime="00:00:52.80" resultid="1540" heatid="2099" lane="4" />
                <RESULT eventid="1235" points="112" swimtime="00:00:58.73" resultid="1541" heatid="2117" lane="5" />
                <RESULT eventid="1254" points="125" swimtime="00:00:45.81" resultid="1542" heatid="2127" lane="3" entrytime="00:00:50.80" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="De Araujo" birthdate="2015-08-09" gender="F" nation="BRA" license="407185" swrid="5725999" athleteid="1570" externalid="407185">
              <RESULTS>
                <RESULT eventid="1213" points="53" swimtime="00:01:06.82" resultid="1571" heatid="2108" lane="6" entrytime="00:01:11.46" entrycourse="SCM" />
                <RESULT eventid="1235" points="63" swimtime="00:01:10.95" resultid="1572" heatid="2118" lane="6" entrytime="00:01:11.85" entrycourse="SCM" />
                <RESULT eventid="1254" points="57" swimtime="00:00:59.25" resultid="1573" heatid="2127" lane="5" entrytime="00:01:00.25" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Corsine Ferreira" birthdate="2010-03-10" gender="F" nation="BRA" license="353591" swrid="5588608" athleteid="1451" externalid="353591">
              <RESULTS>
                <RESULT eventid="1150" points="323" swimtime="00:00:41.31" resultid="1452" heatid="2083" lane="3" entrytime="00:00:40.13" entrycourse="SCM" />
                <RESULT eventid="1196" points="341" swimtime="00:01:29.18" resultid="1453" heatid="2102" lane="5" entrytime="00:01:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Da Cateburcio" birthdate="2004-01-18" gender="F" nation="BRA" license="407186" swrid="5737919" athleteid="1574" externalid="407186">
              <RESULTS>
                <RESULT eventid="1083" points="75" swimtime="00:01:58.78" resultid="1575" heatid="2050" lane="5" entrytime="00:02:04.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1150" status="DSQ" swimtime="00:01:42.66" resultid="1576" heatid="2082" lane="3" />
                <RESULT eventid="1260" points="85" swimtime="00:00:52.12" resultid="1577" heatid="2131" lane="4" entrytime="00:00:54.06" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Marques Picolo Vinha" birthdate="2010-07-01" gender="M" nation="BRA" license="366990" swrid="5603869" athleteid="1503" externalid="366990">
              <RESULTS>
                <RESULT eventid="1091" points="329" swimtime="00:01:04.95" resultid="1504" heatid="2055" lane="6" entrytime="00:01:04.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="299" swimtime="00:05:17.40" resultid="1505" heatid="2096" lane="5" entrytime="00:05:07.02" entrycourse="SCM" />
                <RESULT eventid="1248" points="240" swimtime="00:01:17.68" resultid="1506" heatid="2124" lane="3" entrytime="00:01:24.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Bessa" birthdate="2003-06-19" gender="M" nation="BRA" license="317841" swrid="5312237" athleteid="1337" externalid="317841">
              <RESULTS>
                <RESULT eventid="1091" points="312" swimtime="00:01:06.05" resultid="1338" heatid="2053" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="545" swimtime="00:00:30.53" resultid="1339" heatid="2086" lane="3" entrytime="00:00:29.77" entrycourse="SCM" />
                <RESULT eventid="1265" points="507" swimtime="00:00:25.28" resultid="1340" heatid="2133" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Forti Francisco" birthdate="2015-07-08" gender="M" nation="BRA" license="392104" swrid="5534395" athleteid="1472" externalid="392104">
              <RESULTS>
                <RESULT eventid="1172" points="110" swimtime="00:01:33.39" resultid="1473" heatid="2091" lane="2" entrytime="00:01:50.67" entrycourse="SCM" />
                <RESULT eventid="1238" points="86" swimtime="00:00:56.39" resultid="1474" heatid="2120" lane="4" entrytime="00:00:57.13" entrycourse="SCM" />
                <RESULT eventid="1257" points="116" swimtime="00:00:41.32" resultid="1475" heatid="2129" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio" lastname="Rafael Padial" birthdate="2014-03-07" gender="M" nation="BRA" license="397331" swrid="5641774" athleteid="1519" externalid="397331">
              <RESULTS>
                <RESULT eventid="1172" points="174" swimtime="00:01:20.17" resultid="1520" heatid="2091" lane="3" entrytime="00:01:23.86" entrycourse="SCM" />
                <RESULT eventid="1216" points="128" swimtime="00:00:43.84" resultid="1521" heatid="2109" lane="3" entrytime="00:00:42.10" entrycourse="SCM" />
                <RESULT eventid="1257" points="172" swimtime="00:00:36.23" resultid="1522" heatid="2130" lane="3" entrytime="00:00:35.06" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Quental De Meireles" birthdate="2008-11-20" gender="M" nation="BRA" license="392103" swrid="5603898" athleteid="1468" externalid="392103">
              <RESULTS>
                <RESULT eventid="1140" points="324" swimtime="00:01:09.50" resultid="1469" heatid="2075" lane="2" entrytime="00:01:08.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1225" points="372" swimtime="00:00:30.24" resultid="1470" heatid="2113" lane="2" />
                <RESULT eventid="1265" points="358" swimtime="00:00:28.38" resultid="1471" heatid="2136" lane="6" entrytime="00:00:28.91" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sara" lastname="Padovin Chiste" birthdate="2015-02-04" gender="F" nation="BRA" license="414849" athleteid="1587" externalid="414849">
              <RESULTS>
                <RESULT eventid="1169" points="92" swimtime="00:01:51.08" resultid="1588" heatid="2089" lane="2" />
                <RESULT eventid="1235" points="96" swimtime="00:01:01.76" resultid="1589" heatid="2117" lane="4" />
                <RESULT eventid="1254" points="78" swimtime="00:00:53.44" resultid="1590" heatid="2126" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Tomazeli" birthdate="2013-02-05" gender="M" nation="BRA" license="392109" swrid="5614097" athleteid="1488" externalid="392109">
              <RESULTS>
                <RESULT eventid="1063" points="154" swimtime="00:03:05.10" resultid="1489" heatid="2041" lane="1" entrytime="00:03:03.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                    <SPLIT distance="100" swimtime="00:01:26.73" />
                    <SPLIT distance="150" swimtime="00:02:14.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="147" swimtime="00:03:27.34" resultid="1490" heatid="2071" lane="2" entrytime="00:03:31.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.34" />
                    <SPLIT distance="100" swimtime="00:01:41.37" />
                    <SPLIT distance="150" swimtime="00:02:40.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="164" swimtime="00:00:36.82" resultid="1491" heatid="2080" lane="5" entrytime="00:00:39.08" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tiago" lastname="Ficher Delmont Pais" birthdate="2010-07-15" gender="M" nation="BRA" license="338533" swrid="5588701" athleteid="1341" externalid="338533">
              <RESULTS>
                <RESULT eventid="1070" points="450" swimtime="00:02:23.04" resultid="1342" heatid="2045" lane="3" entrytime="00:02:23.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.89" />
                    <SPLIT distance="100" swimtime="00:01:05.19" />
                    <SPLIT distance="150" swimtime="00:01:50.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="451" swimtime="00:04:36.75" resultid="1343" heatid="2096" lane="3" entrytime="00:04:45.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                    <SPLIT distance="100" swimtime="00:01:03.73" />
                    <SPLIT distance="150" swimtime="00:01:38.94" />
                    <SPLIT distance="200" swimtime="00:02:14.18" />
                    <SPLIT distance="250" swimtime="00:02:49.33" />
                    <SPLIT distance="300" swimtime="00:03:26.09" />
                    <SPLIT distance="350" swimtime="00:04:04.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Henrique Goes" birthdate="2008-10-26" gender="M" nation="BRA" license="392105" swrid="5603853" athleteid="1476" externalid="392105">
              <RESULTS>
                <RESULT eventid="1070" points="260" swimtime="00:02:51.63" resultid="1477" heatid="2043" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                    <SPLIT distance="100" swimtime="00:01:21.18" />
                    <SPLIT distance="150" swimtime="00:02:10.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="218" swimtime="00:00:41.45" resultid="1478" heatid="2085" lane="4" />
                <RESULT eventid="1180" points="284" swimtime="00:05:22.85" resultid="1479" heatid="2095" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                    <SPLIT distance="100" swimtime="00:01:14.32" />
                    <SPLIT distance="150" swimtime="00:01:55.81" />
                    <SPLIT distance="200" swimtime="00:02:37.86" />
                    <SPLIT distance="250" swimtime="00:03:19.86" />
                    <SPLIT distance="300" swimtime="00:04:01.14" />
                    <SPLIT distance="350" swimtime="00:04:42.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Garcia Cavalcante" birthdate="2008-08-11" gender="M" nation="BRA" license="369676" swrid="5603841" athleteid="1349" externalid="369676">
              <RESULTS>
                <RESULT eventid="1091" points="400" swimtime="00:01:00.81" resultid="1350" heatid="2053" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="417" swimtime="00:04:43.91" resultid="1351" heatid="2094" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                    <SPLIT distance="100" swimtime="00:01:05.27" />
                    <SPLIT distance="150" swimtime="00:01:41.18" />
                    <SPLIT distance="200" swimtime="00:02:17.69" />
                    <SPLIT distance="250" swimtime="00:02:54.35" />
                    <SPLIT distance="300" swimtime="00:03:31.15" />
                    <SPLIT distance="350" swimtime="00:04:07.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="373" swimtime="00:01:16.75" resultid="1352" heatid="2104" lane="2" entrytime="00:01:13.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="De Correa" birthdate="2014-12-03" gender="M" nation="BRA" license="403387" swrid="5676286" athleteid="1535" externalid="403387">
              <RESULTS>
                <RESULT eventid="1216" points="109" swimtime="00:00:46.16" resultid="1536" heatid="2109" lane="4" entrytime="00:00:49.76" entrycourse="SCM" />
                <RESULT eventid="1238" points="86" swimtime="00:00:56.43" resultid="1537" heatid="2119" lane="2" entrytime="00:01:02.81" entrycourse="SCM" />
                <RESULT eventid="1257" points="134" swimtime="00:00:39.33" resultid="1538" heatid="2130" lane="4" entrytime="00:00:40.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Diogo" lastname="Sanchez" birthdate="2012-11-29" gender="M" nation="BRA" license="370658" swrid="5603906" athleteid="1356" externalid="370658">
              <RESULTS>
                <RESULT eventid="1063" points="143" swimtime="00:03:09.64" resultid="1357" heatid="2040" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.73" />
                    <SPLIT distance="100" swimtime="00:01:32.49" />
                    <SPLIT distance="150" swimtime="00:02:22.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="121" swimtime="00:00:44.69" resultid="1358" heatid="2059" lane="1" />
                <RESULT eventid="1131" points="136" swimtime="00:03:32.97" resultid="1359" heatid="2071" lane="5" entrytime="00:03:41.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.17" />
                    <SPLIT distance="100" swimtime="00:01:46.54" />
                    <SPLIT distance="150" swimtime="00:02:44.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Mochiutti Carneiro" birthdate="2010-04-22" gender="F" nation="BRA" license="370670" swrid="5588817" athleteid="1454" externalid="370670">
              <RESULTS>
                <RESULT eventid="1134" points="418" swimtime="00:01:12.26" resultid="1455" heatid="2073" lane="4" entrytime="00:01:12.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="421" swimtime="00:05:08.52" resultid="1456" heatid="2093" lane="4" entrytime="00:05:11.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                    <SPLIT distance="100" swimtime="00:01:11.92" />
                    <SPLIT distance="150" swimtime="00:01:49.41" />
                    <SPLIT distance="200" swimtime="00:02:27.56" />
                    <SPLIT distance="250" swimtime="00:03:06.50" />
                    <SPLIT distance="300" swimtime="00:03:46.13" />
                    <SPLIT distance="350" swimtime="00:04:27.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1260" points="476" swimtime="00:00:29.36" resultid="1457" heatid="2132" lane="2" entrytime="00:00:30.44" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolas" lastname="Baldo De França" birthdate="2014-04-21" gender="M" nation="BRA" license="393773" swrid="5507467" athleteid="1507" externalid="393773">
              <RESULTS>
                <RESULT eventid="1172" points="90" swimtime="00:01:39.96" resultid="1508" heatid="2090" lane="4" />
                <RESULT eventid="1193" points="83" swimtime="00:00:49.76" resultid="1509" heatid="2101" lane="4" entrytime="00:00:48.49" entrycourse="SCM" />
                <RESULT eventid="1238" points="79" swimtime="00:00:58.02" resultid="1510" heatid="2120" lane="5" entrytime="00:00:58.84" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
