<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.80519">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Colombo/Maringá" name="Campeonato Superparanaense 2024" course="SCM" deadline="2024-12-03" entrystartdate="2024-11-25" entrytype="INVITATION" hostclub="Swim Time Brasil" hostclub.url="https://www.swimtimebrasil.com/" number="38330" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/newInterface/eventos/38330" startmethod="1" timing="AUTOMATIC" touchpad="ONESIDE" masters="F" withdrawuntil="2024-12-05" state="PR" nation="BRA" hytek.courseorder="S">
      <AGEDATE value="2024-12-07" type="YEAR" />
      <POOL name="Santa Mônica Clube de Campo/Universidade Estadual de Maringá" lanemin="1" lanemax="6" />
      <FACILITY city="Colombo/Maringá" name="Santa Mônica Clube de Campo/Universidade Estadual de Maringá" nation="BRA" state="PR" street="5000, Rodovia Régis Bittencourt/Avenida Colombo, 5790" street2="Mauá/Zona 7" zip="83413-663/87020-900" />
      <POINTTABLE pointtableid="3017" name="AQUA Point Scoring" version="2024" />
      <FEES>
        <FEE currency="BRL" type="ATHLETE" value="10000" />
      </FEES>
      <QUALIFY from="2023-12-07" until="2024-12-06" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99252-0598" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99252-0598" street="Avenida do Batel, 1230" street2="Sala 202" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2024-12-07" daytime="08:10" endtime="03:27" number="1" officialmeeting="07:30" warmupfrom="07:30" warmupuntil="08:00">
          <EVENTS>
            <EVENT eventid="1061" gender="F" number="1" order="1" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4261" agemax="9" agemin="9" name="[Colombo] Mirim 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2824" />
                    <RANKING order="2" place="2" resultid="2789" />
                    <RANKING order="3" place="3" resultid="3745" />
                    <RANKING order="4" place="4" resultid="2845" />
                    <RANKING order="5" place="5" resultid="3752" />
                    <RANKING order="6" place="6" resultid="2761" />
                    <RANKING order="7" place="7" resultid="1392" />
                    <RANKING order="8" place="8" resultid="1892" />
                    <RANKING order="9" place="9" resultid="2901" />
                    <RANKING order="10" place="10" resultid="3041" />
                    <RANKING order="11" place="-1" resultid="2754" />
                    <RANKING order="12" place="-1" resultid="2775" />
                    <RANKING order="13" place="-1" resultid="2810" />
                    <RANKING order="14" place="-1" resultid="2838" />
                    <RANKING order="15" place="-1" resultid="2852" />
                    <RANKING order="16" place="-1" resultid="2915" />
                    <RANKING order="17" place="-1" resultid="2936" />
                    <RANKING order="18" place="-1" resultid="2978" />
                    <RANKING order="19" place="-1" resultid="3005" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5261" agemax="10" agemin="10" name="[Colombo] Mirim 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2567" />
                    <RANKING order="2" place="2" resultid="4058" />
                    <RANKING order="3" place="3" resultid="3928" />
                    <RANKING order="4" place="4" resultid="2859" />
                    <RANKING order="5" place="5" resultid="4167" />
                    <RANKING order="6" place="6" resultid="2574" />
                    <RANKING order="7" place="7" resultid="2670" />
                    <RANKING order="8" place="8" resultid="2719" />
                    <RANKING order="9" place="9" resultid="2796" />
                    <RANKING order="10" place="10" resultid="2677" />
                    <RANKING order="11" place="11" resultid="4208" />
                    <RANKING order="12" place="12" resultid="2095" />
                    <RANKING order="13" place="13" resultid="4065" />
                    <RANKING order="14" place="14" resultid="4153" />
                    <RANKING order="15" place="15" resultid="1398" />
                    <RANKING order="16" place="16" resultid="2733" />
                    <RANKING order="17" place="17" resultid="2740" />
                    <RANKING order="18" place="18" resultid="3421" />
                    <RANKING order="19" place="19" resultid="3759" />
                    <RANKING order="20" place="-1" resultid="2637" />
                    <RANKING order="21" place="-1" resultid="2698" />
                    <RANKING order="22" place="-1" resultid="2998" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4458" agemax="9" agemin="9" name="[Maringá] Mirim 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3296" />
                    <RANKING order="2" place="2" resultid="1735" />
                    <RANKING order="3" place="3" resultid="1704" />
                    <RANKING order="4" place="-1" resultid="1773" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5262" agemax="10" agemin="10" name="[Maringá] Mirim 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3226" />
                    <RANKING order="2" place="2" resultid="1723" />
                    <RANKING order="3" place="3" resultid="1613" />
                    <RANKING order="4" place="4" resultid="1998" />
                    <RANKING order="5" place="5" resultid="1716" />
                    <RANKING order="6" place="6" resultid="3445" />
                    <RANKING order="7" place="7" resultid="3554" />
                    <RANKING order="8" place="8" resultid="3390" />
                    <RANKING order="9" place="9" resultid="3254" />
                    <RANKING order="10" place="10" resultid="3600" />
                    <RANKING order="11" place="-1" resultid="1730" />
                    <RANKING order="12" place="-1" resultid="3472" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4645" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4646" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4647" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4648" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4649" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4650" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4651" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4652" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4653" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4654" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1064" gender="F" number="2" order="2" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5275" agemax="11" agemin="11" name="[Colombo] Petiz 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2964" />
                    <RANKING order="2" place="2" resultid="3955" />
                    <RANKING order="3" place="3" resultid="4238" />
                    <RANKING order="4" place="4" resultid="2462" />
                    <RANKING order="5" place="5" resultid="3275" />
                    <RANKING order="6" place="6" resultid="2441" />
                    <RANKING order="7" place="7" resultid="2434" />
                    <RANKING order="8" place="8" resultid="2483" />
                    <RANKING order="9" place="9" resultid="2546" />
                    <RANKING order="10" place="10" resultid="3935" />
                    <RANKING order="11" place="11" resultid="2644" />
                    <RANKING order="12" place="12" resultid="1851" />
                    <RANKING order="13" place="13" resultid="2497" />
                    <RANKING order="14" place="14" resultid="2047" />
                    <RANKING order="15" place="15" resultid="3696" />
                    <RANKING order="16" place="16" resultid="3976" />
                    <RANKING order="17" place="17" resultid="4003" />
                    <RANKING order="18" place="18" resultid="3363" />
                    <RANKING order="19" place="19" resultid="2712" />
                    <RANKING order="20" place="20" resultid="2616" />
                    <RANKING order="21" place="-1" resultid="3376" />
                    <RANKING order="22" place="-1" resultid="4052" />
                    <RANKING order="23" place="-1" resultid="4181" />
                    <RANKING order="24" place="-1" resultid="1906" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5276" agemax="12" agemin="12" name="[Colombo] Petiz 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2511" />
                    <RANKING order="2" place="2" resultid="2385" />
                    <RANKING order="3" place="3" resultid="2331" />
                    <RANKING order="4" place="4" resultid="4107" />
                    <RANKING order="5" place="5" resultid="2324" />
                    <RANKING order="6" place="6" resultid="2378" />
                    <RANKING order="7" place="7" resultid="1846" />
                    <RANKING order="8" place="8" resultid="2469" />
                    <RANKING order="9" place="9" resultid="3921" />
                    <RANKING order="10" place="10" resultid="2371" />
                    <RANKING order="11" place="11" resultid="2705" />
                    <RANKING order="12" place="12" resultid="2943" />
                    <RANKING order="13" place="13" resultid="2455" />
                    <RANKING order="14" place="13" resultid="3948" />
                    <RANKING order="15" place="15" resultid="3459" />
                    <RANKING order="16" place="16" resultid="2077" />
                    <RANKING order="17" place="17" resultid="2406" />
                    <RANKING order="18" place="18" resultid="3349" />
                    <RANKING order="19" place="19" resultid="3780" />
                    <RANKING order="20" place="20" resultid="1878" />
                    <RANKING order="21" place="21" resultid="1371" />
                    <RANKING order="22" place="22" resultid="4140" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5279" agemax="13" agemin="13" name="[Colombo] Infantil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2282" />
                    <RANKING order="2" place="2" resultid="3149" />
                    <RANKING order="3" place="3" resultid="2873" />
                    <RANKING order="4" place="4" resultid="2303" />
                    <RANKING order="5" place="5" resultid="1385" />
                    <RANKING order="6" place="6" resultid="2448" />
                    <RANKING order="7" place="7" resultid="2254" />
                    <RANKING order="8" place="8" resultid="2866" />
                    <RANKING order="9" place="9" resultid="2275" />
                    <RANKING order="10" place="10" resultid="2268" />
                    <RANKING order="11" place="11" resultid="2154" />
                    <RANKING order="12" place="12" resultid="4160" />
                    <RANKING order="13" place="-1" resultid="1899" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5280" agemax="14" agemin="14" name="[Colombo] Infantil 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2602" />
                    <RANKING order="2" place="2" resultid="3724" />
                    <RANKING order="3" place="3" resultid="2198" />
                    <RANKING order="4" place="4" resultid="2191" />
                    <RANKING order="5" place="5" resultid="4187" />
                    <RANKING order="6" place="6" resultid="3610" />
                    <RANKING order="7" place="7" resultid="4194" />
                    <RANKING order="8" place="8" resultid="1807" />
                    <RANKING order="9" place="9" resultid="3407" />
                    <RANKING order="10" place="10" resultid="3717" />
                    <RANKING order="11" place="-1" resultid="3643" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5281" agemax="15" agemin="15" name="[Colombo] Juvenil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3802" />
                    <RANKING order="2" place="2" resultid="1350" />
                    <RANKING order="3" place="3" resultid="3100" />
                    <RANKING order="4" place="4" resultid="3841" />
                    <RANKING order="5" place="5" resultid="2005" />
                    <RANKING order="6" place="6" resultid="2042" />
                    <RANKING order="7" place="7" resultid="1357" />
                    <RANKING order="8" place="8" resultid="2036" />
                    <RANKING order="9" place="9" resultid="3861" />
                    <RANKING order="10" place="10" resultid="2140" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5282" agemax="-1" agemin="16" name="[Colombo] Juvenil 2/Sênior">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5255" />
                    <RANKING order="2" place="2" resultid="3738" />
                    <RANKING order="3" place="3" resultid="1820" />
                    <RANKING order="4" place="4" resultid="3356" />
                    <RANKING order="5" place="5" resultid="3731" />
                    <RANKING order="6" place="6" resultid="3650" />
                    <RANKING order="7" place="7" resultid="4252" />
                    <RANKING order="8" place="8" resultid="3662" />
                    <RANKING order="9" place="9" resultid="1839" />
                    <RANKING order="10" place="10" resultid="2065" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5283" agemax="11" agemin="11" name="[Maringá] Petiz 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3310" />
                    <RANKING order="2" place="2" resultid="1676" />
                    <RANKING order="3" place="3" resultid="3261" />
                    <RANKING order="4" place="4" resultid="3247" />
                    <RANKING order="5" place="5" resultid="3240" />
                    <RANKING order="6" place="6" resultid="3212" />
                    <RANKING order="7" place="7" resultid="3128" />
                    <RANKING order="8" place="8" resultid="1566" />
                    <RANKING order="9" place="9" resultid="1606" />
                    <RANKING order="10" place="-1" resultid="3486" />
                    <RANKING order="11" place="-1" resultid="1545" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5284" agemax="12" agemin="12" name="[Maringá] Petiz 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3142" />
                    <RANKING order="2" place="2" resultid="3114" />
                    <RANKING order="3" place="3" resultid="3547" />
                    <RANKING order="4" place="4" resultid="1559" />
                    <RANKING order="5" place="5" resultid="1599" />
                    <RANKING order="6" place="6" resultid="3205" />
                    <RANKING order="7" place="7" resultid="3414" />
                    <RANKING order="8" place="8" resultid="3233" />
                    <RANKING order="9" place="9" resultid="3303" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5285" agemax="13" agemin="13" name="[Maringá] Infantil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1496" />
                    <RANKING order="2" place="2" resultid="1489" />
                    <RANKING order="3" place="3" resultid="3282" />
                    <RANKING order="4" place="4" resultid="1972" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5286" agemax="14" agemin="14" name="[Maringá] Infantil 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1932" />
                    <RANKING order="2" place="2" resultid="1482" />
                    <RANKING order="3" place="3" resultid="1959" />
                    <RANKING order="4" place="4" resultid="3177" />
                    <RANKING order="5" place="5" resultid="3568" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5287" agemax="15" agemin="15" name="[Maringá] Juvenil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1952" />
                    <RANKING order="2" place="2" resultid="1517" />
                    <RANKING order="3" place="-1" resultid="1524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5288" agemax="-1" agemin="16" name="[Maringá] Juvenil 2/Sênior">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1510" />
                    <RANKING order="2" place="2" resultid="1945" />
                    <RANKING order="3" place="3" resultid="3521" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4657" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4658" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4659" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4660" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4661" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4662" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4663" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4664" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4665" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4666" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4667" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4668" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="4669" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="4670" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="4671" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="4672" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="4673" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="4674" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="4675" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="4676" number="20" order="20" status="OFFICIAL" />
                <HEAT heatid="4677" number="21" order="21" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="4411" gender="F" number="2" order="3" round="SEM" preveventid="1064">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4412" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5608" />
                    <RANKING order="2" place="2" resultid="5381" />
                    <RANKING order="3" place="3" resultid="5382" />
                    <RANKING order="4" place="4" resultid="5383" />
                    <RANKING order="5" place="5" resultid="5385" />
                    <RANKING order="6" place="6" resultid="5607" />
                    <RANKING order="7" place="7" resultid="5610" />
                    <RANKING order="8" place="8" resultid="5609" />
                    <RANKING order="9" place="9" resultid="5384" />
                    <RANKING order="10" place="10" resultid="5386" />
                    <RANKING order="11" place="11" resultid="5611" />
                    <RANKING order="12" place="12" resultid="5612" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4474" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5387" />
                    <RANKING order="2" place="2" resultid="5388" />
                    <RANKING order="3" place="3" resultid="5389" />
                    <RANKING order="4" place="4" resultid="5614" />
                    <RANKING order="5" place="5" resultid="5613" />
                    <RANKING order="6" place="6" resultid="5390" />
                    <RANKING order="7" place="7" resultid="5392" />
                    <RANKING order="8" place="8" resultid="5391" />
                    <RANKING order="9" place="9" resultid="5616" />
                    <RANKING order="10" place="10" resultid="5615" />
                    <RANKING order="11" place="11" resultid="5618" />
                    <RANKING order="12" place="12" resultid="5617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4476" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5353" />
                    <RANKING order="2" place="2" resultid="5354" />
                    <RANKING order="3" place="3" resultid="5356" />
                    <RANKING order="4" place="4" resultid="5357" />
                    <RANKING order="5" place="5" resultid="5355" />
                    <RANKING order="6" place="6" resultid="5358" />
                    <RANKING order="7" place="7" resultid="5619" />
                    <RANKING order="8" place="8" resultid="5620" />
                    <RANKING order="9" place="9" resultid="5622" />
                    <RANKING order="10" place="10" resultid="5621" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4477" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5624" />
                    <RANKING order="2" place="2" resultid="5623" />
                    <RANKING order="3" place="3" resultid="5625" />
                    <RANKING order="4" place="4" resultid="5326" />
                    <RANKING order="5" place="5" resultid="5328" />
                    <RANKING order="6" place="6" resultid="5327" />
                    <RANKING order="7" place="7" resultid="5329" />
                    <RANKING order="8" place="8" resultid="5330" />
                    <RANKING order="9" place="9" resultid="5331" />
                    <RANKING order="10" place="10" resultid="5626" />
                    <RANKING order="11" place="11" resultid="5627" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4478" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5335" />
                    <RANKING order="2" place="2" resultid="5336" />
                    <RANKING order="3" place="3" resultid="5337" />
                    <RANKING order="4" place="4" resultid="5338" />
                    <RANKING order="5" place="5" resultid="5340" />
                    <RANKING order="6" place="6" resultid="5339" />
                    <RANKING order="7" place="7" resultid="5628" />
                    <RANKING order="8" place="8" resultid="5629" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4479" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5344" />
                    <RANKING order="2" place="2" resultid="5630" />
                    <RANKING order="3" place="3" resultid="5345" />
                    <RANKING order="4" place="4" resultid="5347" />
                    <RANKING order="5" place="5" resultid="5348" />
                    <RANKING order="6" place="6" resultid="5349" />
                    <RANKING order="7" place="7" resultid="5631" />
                    <RANKING order="8" place="8" resultid="5632" />
                    <RANKING order="9" place="-1" resultid="5346" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4678" agegroupid="4412" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4679" agegroupid="4412" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4680" agegroupid="4474" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4681" agegroupid="4474" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4682" agegroupid="4476" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4683" agegroupid="4476" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4684" agegroupid="4477" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4685" agegroupid="4477" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4686" agegroupid="4478" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4687" agegroupid="4478" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4688" agegroupid="4479" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4689" agegroupid="4479" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="4409" gender="F" number="1" order="4" round="FIN" preveventid="1061">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4410" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5365" />
                    <RANKING order="2" place="2" resultid="5364" />
                    <RANKING order="3" place="3" resultid="5363" />
                    <RANKING order="4" place="4" resultid="5366" />
                    <RANKING order="5" place="5" resultid="5368" />
                    <RANKING order="6" place="6" resultid="5367" />
                    <RANKING order="7" place="7" resultid="9015" />
                    <RANKING order="8" place="8" resultid="9016" />
                    <RANKING order="9" place="9" resultid="9017" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4459" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9018" />
                    <RANKING order="2" place="2" resultid="5371" />
                    <RANKING order="3" place="3" resultid="5372" />
                    <RANKING order="4" place="4" resultid="5370" />
                    <RANKING order="5" place="5" resultid="10323" />
                    <RANKING order="6" place="6" resultid="5374" />
                    <RANKING order="7" place="7" resultid="9019" />
                    <RANKING order="8" place="8" resultid="5373" />
                    <RANKING order="9" place="9" resultid="9020" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4655" agegroupid="4410" final="F1" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9001" agegroupid="4410" final="F2" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4656" agegroupid="4459" final="F1" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9002" agegroupid="4459" final="F2" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="4413" gender="F" number="2" order="5" round="FIN" preveventid="4411">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4522" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5633" />
                    <RANKING order="2" place="2" resultid="5634" />
                    <RANKING order="3" place="3" resultid="5376" />
                    <RANKING order="4" place="4" resultid="5635" />
                    <RANKING order="5" place="5" resultid="5377" />
                    <RANKING order="6" place="6" resultid="5375" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4523" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5393" />
                    <RANKING order="2" place="2" resultid="5637" />
                    <RANKING order="3" place="3" resultid="5636" />
                    <RANKING order="4" place="4" resultid="5394" />
                    <RANKING order="5" place="5" resultid="5395" />
                    <RANKING order="6" place="6" resultid="5638" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4524" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5359" />
                    <RANKING order="2" place="2" resultid="5361" />
                    <RANKING order="3" place="3" resultid="5639" />
                    <RANKING order="4" place="4" resultid="5360" />
                    <RANKING order="5" place="5" resultid="5640" />
                    <RANKING order="6" place="6" resultid="5641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4525" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5643" />
                    <RANKING order="2" place="2" resultid="5642" />
                    <RANKING order="3" place="3" resultid="5644" />
                    <RANKING order="4" place="4" resultid="5334" />
                    <RANKING order="5" place="5" resultid="5332" />
                    <RANKING order="6" place="6" resultid="5333" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4526" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5341" />
                    <RANKING order="2" place="2" resultid="5342" />
                    <RANKING order="3" place="3" resultid="5343" />
                    <RANKING order="4" place="4" resultid="5645" />
                    <RANKING order="5" place="5" resultid="5646" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4527" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5647" />
                    <RANKING order="2" place="2" resultid="5350" />
                    <RANKING order="3" place="3" resultid="5351" />
                    <RANKING order="4" place="4" resultid="5648" />
                    <RANKING order="5" place="5" resultid="10322" />
                    <RANKING order="6" place="6" resultid="5649" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4690" agegroupid="4522" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4691" agegroupid="4523" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4692" agegroupid="4524" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4693" agegroupid="4525" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4694" agegroupid="4526" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4695" agegroupid="4527" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1074" gender="F" number="3" order="6" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5263" agemax="9" agemin="9" name="[Colombo] Mirim 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3746" />
                    <RANKING order="2" place="2" resultid="2846" />
                    <RANKING order="3" place="3" resultid="2825" />
                    <RANKING order="4" place="4" resultid="3753" />
                    <RANKING order="5" place="5" resultid="2790" />
                    <RANKING order="6" place="6" resultid="1393" />
                    <RANKING order="7" place="7" resultid="3042" />
                    <RANKING order="8" place="8" resultid="2762" />
                    <RANKING order="9" place="9" resultid="2902" />
                    <RANKING order="10" place="10" resultid="1893" />
                    <RANKING order="11" place="11" resultid="2755" />
                    <RANKING order="12" place="12" resultid="2776" />
                    <RANKING order="13" place="-1" resultid="2811" />
                    <RANKING order="14" place="-1" resultid="2839" />
                    <RANKING order="15" place="-1" resultid="2853" />
                    <RANKING order="16" place="-1" resultid="2916" />
                    <RANKING order="17" place="-1" resultid="2937" />
                    <RANKING order="18" place="-1" resultid="2979" />
                    <RANKING order="19" place="-1" resultid="3006" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5264" agemax="10" agemin="10" name="[Colombo] Mirim 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2568" />
                    <RANKING order="2" place="2" resultid="4059" />
                    <RANKING order="3" place="3" resultid="3929" />
                    <RANKING order="4" place="4" resultid="2797" />
                    <RANKING order="5" place="5" resultid="4168" />
                    <RANKING order="6" place="6" resultid="2860" />
                    <RANKING order="7" place="7" resultid="4066" />
                    <RANKING order="8" place="8" resultid="2575" />
                    <RANKING order="9" place="9" resultid="4209" />
                    <RANKING order="10" place="10" resultid="2671" />
                    <RANKING order="11" place="11" resultid="2720" />
                    <RANKING order="12" place="12" resultid="2678" />
                    <RANKING order="13" place="13" resultid="2741" />
                    <RANKING order="14" place="14" resultid="2734" />
                    <RANKING order="15" place="15" resultid="3422" />
                    <RANKING order="16" place="16" resultid="1399" />
                    <RANKING order="17" place="17" resultid="3760" />
                    <RANKING order="18" place="18" resultid="2096" />
                    <RANKING order="19" place="19" resultid="4154" />
                    <RANKING order="20" place="-1" resultid="2638" />
                    <RANKING order="21" place="-1" resultid="2699" />
                    <RANKING order="22" place="-1" resultid="2999" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5265" agemax="9" agemin="9" name="[Maringá] Mirim 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3297" />
                    <RANKING order="2" place="2" resultid="1705" />
                    <RANKING order="3" place="3" resultid="1736" />
                    <RANKING order="4" place="-1" resultid="1774" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5266" agemax="10" agemin="10" name="[Maringá] Mirim 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1724" />
                    <RANKING order="2" place="2" resultid="3227" />
                    <RANKING order="3" place="3" resultid="3255" />
                    <RANKING order="4" place="4" resultid="1999" />
                    <RANKING order="5" place="5" resultid="3555" />
                    <RANKING order="6" place="6" resultid="1614" />
                    <RANKING order="7" place="7" resultid="3601" />
                    <RANKING order="8" place="8" resultid="3446" />
                    <RANKING order="9" place="9" resultid="1717" />
                    <RANKING order="10" place="10" resultid="3391" />
                    <RANKING order="11" place="-1" resultid="3473" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4696" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4697" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4698" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4699" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4700" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4701" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4702" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4703" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4704" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4705" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1077" gender="F" number="4" order="7" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5289" agemax="11" agemin="11" name="[Colombo] Petiz 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2484" />
                    <RANKING order="2" place="2" resultid="2547" />
                    <RANKING order="3" place="3" resultid="2435" />
                    <RANKING order="4" place="4" resultid="2498" />
                    <RANKING order="5" place="5" resultid="3956" />
                    <RANKING order="6" place="6" resultid="3276" />
                    <RANKING order="7" place="7" resultid="2463" />
                    <RANKING order="8" place="8" resultid="3936" />
                    <RANKING order="9" place="9" resultid="3377" />
                    <RANKING order="10" place="10" resultid="2442" />
                    <RANKING order="11" place="11" resultid="2965" />
                    <RANKING order="12" place="12" resultid="2048" />
                    <RANKING order="13" place="13" resultid="1852" />
                    <RANKING order="14" place="14" resultid="3977" />
                    <RANKING order="15" place="15" resultid="4004" />
                    <RANKING order="16" place="16" resultid="4239" />
                    <RANKING order="17" place="17" resultid="3697" />
                    <RANKING order="18" place="18" resultid="3364" />
                    <RANKING order="19" place="19" resultid="2645" />
                    <RANKING order="20" place="20" resultid="2617" />
                    <RANKING order="21" place="21" resultid="1907" />
                    <RANKING order="22" place="22" resultid="2713" />
                    <RANKING order="23" place="23" resultid="4182" />
                    <RANKING order="24" place="24" resultid="4053" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5290" agemax="12" agemin="12" name="[Colombo] Petiz 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2512" />
                    <RANKING order="2" place="2" resultid="2332" />
                    <RANKING order="3" place="3" resultid="2706" />
                    <RANKING order="4" place="4" resultid="2470" />
                    <RANKING order="5" place="5" resultid="2325" />
                    <RANKING order="6" place="6" resultid="4108" />
                    <RANKING order="7" place="7" resultid="2386" />
                    <RANKING order="8" place="8" resultid="3949" />
                    <RANKING order="9" place="9" resultid="2407" />
                    <RANKING order="10" place="10" resultid="2456" />
                    <RANKING order="11" place="11" resultid="2379" />
                    <RANKING order="12" place="12" resultid="1847" />
                    <RANKING order="13" place="13" resultid="3922" />
                    <RANKING order="14" place="14" resultid="2944" />
                    <RANKING order="15" place="15" resultid="3460" />
                    <RANKING order="16" place="16" resultid="2078" />
                    <RANKING order="17" place="17" resultid="2372" />
                    <RANKING order="18" place="18" resultid="1879" />
                    <RANKING order="19" place="19" resultid="3781" />
                    <RANKING order="20" place="20" resultid="3350" />
                    <RANKING order="21" place="21" resultid="1372" />
                    <RANKING order="22" place="22" resultid="4141" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5291" agemax="13" agemin="13" name="[Colombo] Infantil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2304" />
                    <RANKING order="2" place="2" resultid="2449" />
                    <RANKING order="3" place="3" resultid="1386" />
                    <RANKING order="4" place="4" resultid="2255" />
                    <RANKING order="5" place="5" resultid="2283" />
                    <RANKING order="6" place="6" resultid="2276" />
                    <RANKING order="7" place="7" resultid="2867" />
                    <RANKING order="8" place="8" resultid="3150" />
                    <RANKING order="9" place="9" resultid="2155" />
                    <RANKING order="10" place="10" resultid="2874" />
                    <RANKING order="11" place="11" resultid="1900" />
                    <RANKING order="12" place="12" resultid="4161" />
                    <RANKING order="13" place="13" resultid="2269" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5292" agemax="14" agemin="14" name="[Colombo] Infantil 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2199" />
                    <RANKING order="2" place="2" resultid="4188" />
                    <RANKING order="3" place="3" resultid="2192" />
                    <RANKING order="4" place="4" resultid="4195" />
                    <RANKING order="5" place="5" resultid="3408" />
                    <RANKING order="6" place="6" resultid="2603" />
                    <RANKING order="7" place="7" resultid="1808" />
                    <RANKING order="8" place="8" resultid="3644" />
                    <RANKING order="9" place="9" resultid="3611" />
                    <RANKING order="10" place="10" resultid="3725" />
                    <RANKING order="11" place="11" resultid="3718" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5293" agemax="15" agemin="15" name="[Colombo] Juvenil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3803" />
                    <RANKING order="2" place="2" resultid="1351" />
                    <RANKING order="3" place="3" resultid="2006" />
                    <RANKING order="4" place="4" resultid="3101" />
                    <RANKING order="5" place="5" resultid="2043" />
                    <RANKING order="6" place="5" resultid="3842" />
                    <RANKING order="7" place="7" resultid="1358" />
                    <RANKING order="8" place="8" resultid="3862" />
                    <RANKING order="9" place="9" resultid="2037" />
                    <RANKING order="10" place="10" resultid="2141" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5294" agemax="-1" agemin="16" name="[Colombo] Juvenil 2/Sênior">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5325" />
                    <RANKING order="2" place="2" resultid="3739" />
                    <RANKING order="3" place="3" resultid="1821" />
                    <RANKING order="4" place="4" resultid="3651" />
                    <RANKING order="5" place="5" resultid="3357" />
                    <RANKING order="6" place="6" resultid="3732" />
                    <RANKING order="7" place="7" resultid="3663" />
                    <RANKING order="8" place="8" resultid="1840" />
                    <RANKING order="9" place="9" resultid="4253" />
                    <RANKING order="10" place="10" resultid="2066" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5295" agemax="11" agemin="11" name="[Maringá] Petiz 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1677" />
                    <RANKING order="2" place="2" resultid="3311" />
                    <RANKING order="3" place="3" resultid="3248" />
                    <RANKING order="4" place="4" resultid="3241" />
                    <RANKING order="5" place="5" resultid="3262" />
                    <RANKING order="6" place="6" resultid="1567" />
                    <RANKING order="7" place="7" resultid="3213" />
                    <RANKING order="8" place="8" resultid="1607" />
                    <RANKING order="9" place="-1" resultid="3129" />
                    <RANKING order="10" place="-1" resultid="3487" />
                    <RANKING order="11" place="-1" resultid="1546" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5296" agemax="12" agemin="12" name="[Maringá] Petiz 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3115" />
                    <RANKING order="2" place="2" resultid="3143" />
                    <RANKING order="3" place="3" resultid="1560" />
                    <RANKING order="4" place="4" resultid="3548" />
                    <RANKING order="5" place="5" resultid="3234" />
                    <RANKING order="6" place="6" resultid="1600" />
                    <RANKING order="7" place="7" resultid="3415" />
                    <RANKING order="8" place="8" resultid="3304" />
                    <RANKING order="9" place="9" resultid="3206" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5297" agemax="13" agemin="13" name="[Maringá] Infantil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1490" />
                    <RANKING order="2" place="2" resultid="3283" />
                    <RANKING order="3" place="3" resultid="1497" />
                    <RANKING order="4" place="4" resultid="1973" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5298" agemax="14" agemin="14" name="[Maringá] Infantil 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1933" />
                    <RANKING order="2" place="2" resultid="1960" />
                    <RANKING order="3" place="3" resultid="1483" />
                    <RANKING order="4" place="4" resultid="3178" />
                    <RANKING order="5" place="5" resultid="3569" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5299" agemax="15" agemin="15" name="[Maringá] Juvenil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1518" />
                    <RANKING order="2" place="2" resultid="1953" />
                    <RANKING order="3" place="-1" resultid="1525" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5300" agemax="-1" agemin="16" name="[Maringá] Juvenil 2/Sênior">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1511" />
                    <RANKING order="2" place="2" resultid="1946" />
                    <RANKING order="3" place="3" resultid="3522" />
                    <RANKING order="4" place="4" resultid="1764" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4708" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4709" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4710" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4711" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4712" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4713" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4714" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4715" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4716" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4717" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4718" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4719" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="4720" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="4721" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="4722" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="4723" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="4724" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="4725" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="4726" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="4727" number="20" order="20" status="OFFICIAL" />
                <HEAT heatid="4728" number="21" order="21" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="4417" gender="F" number="4" order="8" round="SEM" preveventid="1077">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4480" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5409" />
                    <RANKING order="2" place="2" resultid="5408" />
                    <RANKING order="3" place="3" resultid="5650" />
                    <RANKING order="4" place="4" resultid="5410" />
                    <RANKING order="5" place="5" resultid="5412" />
                    <RANKING order="6" place="6" resultid="5652" />
                    <RANKING order="7" place="7" resultid="5651" />
                    <RANKING order="8" place="8" resultid="5413" />
                    <RANKING order="9" place="9" resultid="5411" />
                    <RANKING order="10" place="10" resultid="5653" />
                    <RANKING order="11" place="11" resultid="5654" />
                    <RANKING order="12" place="12" resultid="5655" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4481" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5417" />
                    <RANKING order="2" place="2" resultid="5418" />
                    <RANKING order="3" place="3" resultid="5421" />
                    <RANKING order="4" place="4" resultid="5419" />
                    <RANKING order="5" place="5" resultid="5656" />
                    <RANKING order="6" place="6" resultid="5420" />
                    <RANKING order="7" place="7" resultid="5422" />
                    <RANKING order="8" place="8" resultid="5657" />
                    <RANKING order="9" place="9" resultid="5658" />
                    <RANKING order="10" place="10" resultid="5659" />
                    <RANKING order="11" place="11" resultid="5661" />
                    <RANKING order="12" place="-1" resultid="5660" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4482" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5426" />
                    <RANKING order="2" place="2" resultid="5432" />
                    <RANKING order="3" place="3" resultid="5428" />
                    <RANKING order="4" place="4" resultid="5429" />
                    <RANKING order="5" place="5" resultid="5430" />
                    <RANKING order="6" place="6" resultid="5431" />
                    <RANKING order="7" place="7" resultid="5664" />
                    <RANKING order="8" place="8" resultid="5662" />
                    <RANKING order="9" place="9" resultid="5663" />
                    <RANKING order="10" place="10" resultid="5665" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4483" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5436" />
                    <RANKING order="2" place="2" resultid="5438" />
                    <RANKING order="3" place="3" resultid="5437" />
                    <RANKING order="4" place="4" resultid="5668" />
                    <RANKING order="5" place="5" resultid="5667" />
                    <RANKING order="6" place="6" resultid="5669" />
                    <RANKING order="7" place="7" resultid="5439" />
                    <RANKING order="8" place="8" resultid="5440" />
                    <RANKING order="9" place="9" resultid="5441" />
                    <RANKING order="10" place="10" resultid="5666" />
                    <RANKING order="11" place="11" resultid="5670" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4484" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5445" />
                    <RANKING order="2" place="2" resultid="5446" />
                    <RANKING order="3" place="3" resultid="5447" />
                    <RANKING order="4" place="4" resultid="5449" />
                    <RANKING order="5" place="5" resultid="5448" />
                    <RANKING order="6" place="6" resultid="5450" />
                    <RANKING order="7" place="7" resultid="5671" />
                    <RANKING order="8" place="8" resultid="5672" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4485" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5454" />
                    <RANKING order="2" place="2" resultid="5458" />
                    <RANKING order="3" place="3" resultid="5455" />
                    <RANKING order="4" place="4" resultid="5456" />
                    <RANKING order="5" place="5" resultid="5457" />
                    <RANKING order="6" place="6" resultid="5673" />
                    <RANKING order="7" place="7" resultid="5459" />
                    <RANKING order="8" place="8" resultid="5674" />
                    <RANKING order="9" place="9" resultid="5675" />
                    <RANKING order="10" place="10" resultid="5676" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4729" agegroupid="4480" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4730" agegroupid="4480" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4731" agegroupid="4481" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4732" agegroupid="4481" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4733" agegroupid="4482" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4734" agegroupid="4482" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4735" agegroupid="4483" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4736" agegroupid="4483" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4737" agegroupid="4484" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4738" agegroupid="4484" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4739" agegroupid="4485" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4740" agegroupid="4485" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="4415" gender="F" number="3" order="9" round="FIN" preveventid="1074">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4460" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5396" />
                    <RANKING order="2" place="2" resultid="5397" />
                    <RANKING order="3" place="3" resultid="5398" />
                    <RANKING order="4" place="4" resultid="5399" />
                    <RANKING order="5" place="5" resultid="5400" />
                    <RANKING order="6" place="6" resultid="5401" />
                    <RANKING order="7" place="7" resultid="9009" />
                    <RANKING order="8" place="8" resultid="9010" />
                    <RANKING order="9" place="9" resultid="9011" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4461" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5402" />
                    <RANKING order="2" place="2" resultid="9013" />
                    <RANKING order="3" place="3" resultid="5403" />
                    <RANKING order="4" place="4" resultid="5404" />
                    <RANKING order="5" place="5" resultid="5406" />
                    <RANKING order="6" place="6" resultid="5407" />
                    <RANKING order="7" place="7" resultid="5405" />
                    <RANKING order="8" place="8" resultid="9012" />
                    <RANKING order="9" place="9" resultid="9021" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4706" agegroupid="4460" final="F1" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9003" agegroupid="4460" final="F2" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4707" agegroupid="4461" final="F1" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9004" agegroupid="4461" final="F2" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="4419" gender="F" number="4" order="10" round="FIN" preveventid="4417">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4528" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5677" />
                    <RANKING order="2" place="2" resultid="5416" />
                    <RANKING order="3" place="3" resultid="5414" />
                    <RANKING order="4" place="4" resultid="5678" />
                    <RANKING order="5" place="5" resultid="5415" />
                    <RANKING order="6" place="6" resultid="5679" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4529" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5423" />
                    <RANKING order="2" place="2" resultid="5424" />
                    <RANKING order="3" place="3" resultid="5425" />
                    <RANKING order="4" place="4" resultid="5680" />
                    <RANKING order="5" place="5" resultid="5681" />
                    <RANKING order="6" place="6" resultid="5682" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4530" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5433" />
                    <RANKING order="2" place="2" resultid="5434" />
                    <RANKING order="3" place="3" resultid="5435" />
                    <RANKING order="4" place="4" resultid="5684" />
                    <RANKING order="5" place="5" resultid="5683" />
                    <RANKING order="6" place="6" resultid="5685" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4531" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5442" />
                    <RANKING order="2" place="2" resultid="5687" />
                    <RANKING order="3" place="3" resultid="5686" />
                    <RANKING order="4" place="4" resultid="5444" />
                    <RANKING order="5" place="5" resultid="5688" />
                    <RANKING order="6" place="6" resultid="5443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4532" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5452" />
                    <RANKING order="2" place="2" resultid="5451" />
                    <RANKING order="3" place="3" resultid="5453" />
                    <RANKING order="4" place="4" resultid="5690" />
                    <RANKING order="5" place="5" resultid="5689" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4533" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5460" />
                    <RANKING order="2" place="2" resultid="5691" />
                    <RANKING order="3" place="3" resultid="5461" />
                    <RANKING order="4" place="4" resultid="5462" />
                    <RANKING order="5" place="5" resultid="5693" />
                    <RANKING order="6" place="6" resultid="5692" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4741" agegroupid="4528" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4742" agegroupid="4529" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4743" agegroupid="4530" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4744" agegroupid="4531" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4745" agegroupid="4532" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4746" agegroupid="4533" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1087" gender="F" number="5" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="8" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1088" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3083" />
                    <RANKING order="2" place="2" resultid="3496" />
                    <RANKING order="3" place="-1" resultid="3079" />
                    <RANKING order="4" place="-1" resultid="4257" />
                    <RANKING order="5" place="-1" resultid="1801" />
                    <RANKING order="6" place="-1" resultid="3492" />
                    <RANKING order="7" place="-1" resultid="1402" />
                    <RANKING order="8" place="-1" resultid="2115" />
                    <RANKING order="9" place="-1" resultid="2119" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4747" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4748" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5247" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1089" gender="M" number="6" order="12" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5267" agemax="9" agemin="9" name="[Colombo] Mirim 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2768" />
                    <RANKING order="2" place="2" resultid="4024" />
                    <RANKING order="3" place="3" resultid="3012" />
                    <RANKING order="4" place="4" resultid="2747" />
                    <RANKING order="5" place="5" resultid="2831" />
                    <RANKING order="6" place="6" resultid="1911" />
                    <RANKING order="7" place="7" resultid="2817" />
                    <RANKING order="8" place="8" resultid="2929" />
                    <RANKING order="9" place="9" resultid="4226" />
                    <RANKING order="10" place="10" resultid="3481" />
                    <RANKING order="11" place="11" resultid="2922" />
                    <RANKING order="12" place="12" resultid="2950" />
                    <RANKING order="13" place="13" resultid="3317" />
                    <RANKING order="14" place="14" resultid="2957" />
                    <RANKING order="15" place="-1" resultid="2887" />
                    <RANKING order="16" place="-1" resultid="2894" />
                    <RANKING order="17" place="-1" resultid="2908" />
                    <RANKING order="18" place="-1" resultid="2971" />
                    <RANKING order="19" place="-1" resultid="2991" />
                    <RANKING order="20" place="-1" resultid="3060" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5268" agemax="10" agemin="10" name="[Colombo] Mirim 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2691" />
                    <RANKING order="2" place="2" resultid="2595" />
                    <RANKING order="3" place="3" resultid="3424" />
                    <RANKING order="4" place="4" resultid="2581" />
                    <RANKING order="5" place="5" resultid="2684" />
                    <RANKING order="6" place="6" resultid="2588" />
                    <RANKING order="7" place="7" resultid="2880" />
                    <RANKING order="8" place="8" resultid="4072" />
                    <RANKING order="9" place="9" resultid="3962" />
                    <RANKING order="10" place="10" resultid="3969" />
                    <RANKING order="11" place="11" resultid="3989" />
                    <RANKING order="12" place="12" resultid="2656" />
                    <RANKING order="13" place="13" resultid="4093" />
                    <RANKING order="14" place="14" resultid="3019" />
                    <RANKING order="15" place="15" resultid="4100" />
                    <RANKING order="16" place="16" resultid="3073" />
                    <RANKING order="17" place="17" resultid="2663" />
                    <RANKING order="18" place="18" resultid="4121" />
                    <RANKING order="19" place="-1" resultid="1872" />
                    <RANKING order="20" place="-1" resultid="2623" />
                    <RANKING order="21" place="-1" resultid="2630" />
                    <RANKING order="22" place="-1" resultid="2649" />
                    <RANKING order="23" place="-1" resultid="2782" />
                    <RANKING order="24" place="-1" resultid="2803" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5269" agemax="9" agemin="9" name="[Maringá] Mirim 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3289" />
                    <RANKING order="2" place="2" resultid="1697" />
                    <RANKING order="3" place="3" resultid="3268" />
                    <RANKING order="4" place="4" resultid="1669" />
                    <RANKING order="5" place="5" resultid="1627" />
                    <RANKING order="6" place="6" resultid="1787" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5270" agemax="10" agemin="10" name="[Maringá] Mirim 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1620" />
                    <RANKING order="2" place="2" resultid="1709" />
                    <RANKING order="3" place="3" resultid="1683" />
                    <RANKING order="4" place="4" resultid="3431" />
                    <RANKING order="5" place="5" resultid="1662" />
                    <RANKING order="6" place="6" resultid="3342" />
                    <RANKING order="7" place="7" resultid="1744" />
                    <RANKING order="8" place="8" resultid="3397" />
                    <RANKING order="9" place="9" resultid="3438" />
                    <RANKING order="10" place="-1" resultid="1780" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4749" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4750" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4751" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4752" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4753" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4754" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4755" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4756" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4757" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4758" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4759" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1092" gender="M" number="7" order="13" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5301" agemax="11" agemin="11" name="[Colombo] Petiz 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1378" />
                    <RANKING order="2" place="2" resultid="2054" />
                    <RANKING order="3" place="3" resultid="2525" />
                    <RANKING order="4" place="4" resultid="4017" />
                    <RANKING order="5" place="5" resultid="2726" />
                    <RANKING order="6" place="6" resultid="2427" />
                    <RANKING order="7" place="7" resultid="2476" />
                    <RANKING order="8" place="8" resultid="2518" />
                    <RANKING order="9" place="9" resultid="2539" />
                    <RANKING order="10" place="10" resultid="3034" />
                    <RANKING order="11" place="11" resultid="3982" />
                    <RANKING order="12" place="12" resultid="3996" />
                    <RANKING order="13" place="13" resultid="4010" />
                    <RANKING order="14" place="14" resultid="2490" />
                    <RANKING order="15" place="15" resultid="3383" />
                    <RANKING order="16" place="16" resultid="2532" />
                    <RANKING order="17" place="17" resultid="4126" />
                    <RANKING order="18" place="18" resultid="3322" />
                    <RANKING order="19" place="19" resultid="3048" />
                    <RANKING order="20" place="-1" resultid="3710" />
                    <RANKING order="21" place="-1" resultid="3465" />
                    <RANKING order="22" place="-1" resultid="3055" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5302" agemax="12" agemin="12" name="[Colombo] Petiz 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2310" />
                    <RANKING order="2" place="2" resultid="2345" />
                    <RANKING order="3" place="3" resultid="2399" />
                    <RANKING order="4" place="4" resultid="1865" />
                    <RANKING order="5" place="5" resultid="2317" />
                    <RANKING order="6" place="6" resultid="3904" />
                    <RANKING order="7" place="7" resultid="2553" />
                    <RANKING order="8" place="8" resultid="3676" />
                    <RANKING order="9" place="9" resultid="1918" />
                    <RANKING order="10" place="10" resultid="2357" />
                    <RANKING order="11" place="11" resultid="3941" />
                    <RANKING order="12" place="12" resultid="2364" />
                    <RANKING order="13" place="13" resultid="2338" />
                    <RANKING order="14" place="14" resultid="1827" />
                    <RANKING order="15" place="15" resultid="2392" />
                    <RANKING order="16" place="16" resultid="4045" />
                    <RANKING order="17" place="17" resultid="1833" />
                    <RANKING order="18" place="18" resultid="2413" />
                    <RANKING order="19" place="19" resultid="5259" />
                    <RANKING order="20" place="20" resultid="2352" />
                    <RANKING order="21" place="21" resultid="2504" />
                    <RANKING order="22" place="-1" resultid="4086" />
                    <RANKING order="23" place="-1" resultid="4147" />
                    <RANKING order="24" place="-1" resultid="4232" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5303" agemax="13" agemin="13" name="[Colombo] Infantil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4114" />
                    <RANKING order="2" place="2" resultid="2420" />
                    <RANKING order="3" place="3" resultid="3868" />
                    <RANKING order="4" place="4" resultid="1858" />
                    <RANKING order="5" place="5" resultid="2247" />
                    <RANKING order="6" place="6" resultid="2240" />
                    <RANKING order="7" place="7" resultid="3911" />
                    <RANKING order="8" place="8" resultid="2233" />
                    <RANKING order="9" place="9" resultid="3882" />
                    <RANKING order="10" place="10" resultid="1885" />
                    <RANKING order="11" place="11" resultid="2168" />
                    <RANKING order="12" place="12" resultid="2161" />
                    <RANKING order="13" place="13" resultid="3889" />
                    <RANKING order="14" place="14" resultid="2059" />
                    <RANKING order="15" place="15" resultid="2024" />
                    <RANKING order="16" place="16" resultid="2289" />
                    <RANKING order="17" place="17" resultid="3914" />
                    <RANKING order="18" place="18" resultid="2296" />
                    <RANKING order="19" place="19" resultid="3766" />
                    <RANKING order="20" place="20" resultid="2261" />
                    <RANKING order="21" place="21" resultid="3369" />
                    <RANKING order="22" place="-1" resultid="2560" />
                    <RANKING order="23" place="-1" resultid="3452" />
                    <RANKING order="24" place="-1" resultid="4133" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5304" agemax="14" agemin="14" name="[Colombo] Infantil 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2609" />
                    <RANKING order="2" place="2" resultid="2226" />
                    <RANKING order="3" place="3" resultid="2184" />
                    <RANKING order="4" place="4" resultid="3896" />
                    <RANKING order="5" place="5" resultid="4215" />
                    <RANKING order="6" place="6" resultid="4031" />
                    <RANKING order="7" place="7" resultid="3773" />
                    <RANKING order="8" place="8" resultid="4245" />
                    <RANKING order="9" place="9" resultid="2212" />
                    <RANKING order="10" place="10" resultid="2100" />
                    <RANKING order="11" place="11" resultid="4079" />
                    <RANKING order="12" place="12" resultid="2106" />
                    <RANKING order="13" place="13" resultid="2205" />
                    <RANKING order="14" place="14" resultid="2072" />
                    <RANKING order="15" place="-1" resultid="2219" />
                    <RANKING order="16" place="-1" resultid="3875" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5305" agemax="15" agemin="15" name="[Colombo] Juvenil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3827" />
                    <RANKING order="2" place="2" resultid="1364" />
                    <RANKING order="3" place="3" resultid="1343" />
                    <RANKING order="4" place="4" resultid="4038" />
                    <RANKING order="5" place="5" resultid="2017" />
                    <RANKING order="6" place="6" resultid="2030" />
                    <RANKING order="7" place="7" resultid="3622" />
                    <RANKING order="8" place="8" resultid="3854" />
                    <RANKING order="9" place="9" resultid="4174" />
                    <RANKING order="10" place="10" resultid="3629" />
                    <RANKING order="11" place="11" resultid="2176" />
                    <RANKING order="12" place="-1" resultid="3834" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5306" agemax="-1" agemin="16" name="[Colombo] Juvenil 2/Sênior">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3901" />
                    <RANKING order="2" place="2" resultid="3617" />
                    <RANKING order="3" place="3" resultid="3689" />
                    <RANKING order="4" place="4" resultid="3815" />
                    <RANKING order="5" place="5" resultid="3847" />
                    <RANKING order="6" place="6" resultid="3703" />
                    <RANKING order="7" place="7" resultid="3335" />
                    <RANKING order="8" place="8" resultid="2010" />
                    <RANKING order="9" place="9" resultid="3636" />
                    <RANKING order="10" place="10" resultid="2133" />
                    <RANKING order="11" place="11" resultid="3787" />
                    <RANKING order="12" place="12" resultid="3669" />
                    <RANKING order="13" place="13" resultid="2147" />
                    <RANKING order="14" place="14" resultid="3328" />
                    <RANKING order="15" place="15" resultid="3794" />
                    <RANKING order="16" place="16" resultid="4201" />
                    <RANKING order="17" place="17" resultid="3683" />
                    <RANKING order="18" place="18" resultid="3657" />
                    <RANKING order="19" place="-1" resultid="2084" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5307" agemax="11" agemin="11" name="[Maringá] Petiz 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1655" />
                    <RANKING order="2" place="2" resultid="1641" />
                    <RANKING order="3" place="3" resultid="1648" />
                    <RANKING order="4" place="4" resultid="1690" />
                    <RANKING order="5" place="5" resultid="1580" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5308" agemax="12" agemin="12" name="[Maringá] Petiz 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1573" />
                    <RANKING order="2" place="2" resultid="1587" />
                    <RANKING order="3" place="3" resultid="1552" />
                    <RANKING order="4" place="4" resultid="3135" />
                    <RANKING order="5" place="5" resultid="1594" />
                    <RANKING order="6" place="6" resultid="3561" />
                    <RANKING order="7" place="7" resultid="3219" />
                    <RANKING order="8" place="8" resultid="1634" />
                    <RANKING order="9" place="9" resultid="3502" />
                    <RANKING order="10" place="10" resultid="1426" />
                    <RANKING order="11" place="11" resultid="3588" />
                    <RANKING order="12" place="-1" resultid="3581" />
                    <RANKING order="13" place="-1" resultid="3594" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5309" agemax="13" agemin="13" name="[Maringá] Infantil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1406" />
                    <RANKING order="2" place="2" resultid="3163" />
                    <RANKING order="3" place="3" resultid="3170" />
                    <RANKING order="4" place="4" resultid="3191" />
                    <RANKING order="5" place="5" resultid="1461" />
                    <RANKING order="6" place="6" resultid="1984" />
                    <RANKING order="7" place="7" resultid="1454" />
                    <RANKING order="8" place="8" resultid="3107" />
                    <RANKING order="9" place="9" resultid="1991" />
                    <RANKING order="10" place="10" resultid="3121" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5310" agemax="14" agemin="14" name="[Maringá] Infantil 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3093" />
                    <RANKING order="2" place="2" resultid="1468" />
                    <RANKING order="3" place="3" resultid="3574" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5311" agemax="15" agemin="15" name="[Maringá] Juvenil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1419" />
                    <RANKING order="2" place="2" resultid="3508" />
                    <RANKING order="3" place="3" resultid="3535" />
                    <RANKING order="4" place="4" resultid="1440" />
                    <RANKING order="5" place="5" resultid="3156" />
                    <RANKING order="6" place="-1" resultid="1538" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5312" agemax="-1" agemin="16" name="[Maringá] Juvenil 2/Sênior">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1939" />
                    <RANKING order="2" place="2" resultid="1926" />
                    <RANKING order="3" place="3" resultid="1966" />
                    <RANKING order="4" place="4" resultid="1503" />
                    <RANKING order="5" place="5" resultid="1433" />
                    <RANKING order="6" place="6" resultid="1978" />
                    <RANKING order="7" place="7" resultid="1531" />
                    <RANKING order="8" place="8" resultid="3198" />
                    <RANKING order="9" place="9" resultid="1413" />
                    <RANKING order="10" place="10" resultid="1475" />
                    <RANKING order="11" place="11" resultid="1447" />
                    <RANKING order="12" place="12" resultid="3184" />
                    <RANKING order="13" place="13" resultid="1757" />
                    <RANKING order="14" place="14" resultid="3542" />
                    <RANKING order="15" place="15" resultid="3528" />
                    <RANKING order="16" place="16" resultid="1751" />
                    <RANKING order="17" place="-1" resultid="3514" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4762" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4763" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4764" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4765" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4766" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4767" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4768" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4769" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4770" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4771" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4772" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4773" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="4774" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="4775" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="4776" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="4777" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="4778" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="4779" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="4780" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="4781" number="20" order="20" status="OFFICIAL" />
                <HEAT heatid="4782" number="21" order="21" status="OFFICIAL" />
                <HEAT heatid="4783" number="22" order="22" status="OFFICIAL" />
                <HEAT heatid="4784" number="23" order="23" status="OFFICIAL" />
                <HEAT heatid="4785" number="24" order="24" status="OFFICIAL" />
                <HEAT heatid="4786" number="25" order="25" status="OFFICIAL" />
                <HEAT heatid="4787" number="26" order="26" status="OFFICIAL" />
                <HEAT heatid="4788" number="27" order="27" status="OFFICIAL" />
                <HEAT heatid="4789" number="28" order="28" status="OFFICIAL" />
                <HEAT heatid="4790" number="29" order="29" status="OFFICIAL" />
                <HEAT heatid="4791" number="30" order="30" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="4423" gender="M" number="7" order="14" round="SEM" preveventid="1092">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4486" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5482" />
                    <RANKING order="2" place="2" resultid="5484" />
                    <RANKING order="3" place="3" resultid="5485" />
                    <RANKING order="4" place="4" resultid="5486" />
                    <RANKING order="5" place="5" resultid="5481" />
                    <RANKING order="6" place="6" resultid="5483" />
                    <RANKING order="7" place="7" resultid="5694" />
                    <RANKING order="8" place="8" resultid="5695" />
                    <RANKING order="9" place="9" resultid="5696" />
                    <RANKING order="10" place="10" resultid="5697" />
                    <RANKING order="11" place="11" resultid="5698" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4487" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5493" />
                    <RANKING order="2" place="2" resultid="5699" />
                    <RANKING order="3" place="3" resultid="5700" />
                    <RANKING order="4" place="4" resultid="5494" />
                    <RANKING order="5" place="5" resultid="10324" />
                    <RANKING order="6" place="6" resultid="5498" />
                    <RANKING order="7" place="7" resultid="5496" />
                    <RANKING order="8" place="8" resultid="5495" />
                    <RANKING order="9" place="9" resultid="5702" />
                    <RANKING order="10" place="10" resultid="5701" />
                    <RANKING order="11" place="11" resultid="5703" />
                    <RANKING order="12" place="12" resultid="5704" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4488" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5529" />
                    <RANKING order="2" place="2" resultid="5531" />
                    <RANKING order="3" place="3" resultid="5530" />
                    <RANKING order="4" place="4" resultid="5532" />
                    <RANKING order="5" place="5" resultid="5706" />
                    <RANKING order="6" place="6" resultid="5533" />
                    <RANKING order="7" place="7" resultid="5707" />
                    <RANKING order="8" place="8" resultid="5705" />
                    <RANKING order="9" place="9" resultid="5709" />
                    <RANKING order="10" place="10" resultid="5534" />
                    <RANKING order="11" place="11" resultid="5712" />
                    <RANKING order="12" place="12" resultid="5710" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4489" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5541" />
                    <RANKING order="2" place="2" resultid="5538" />
                    <RANKING order="3" place="3" resultid="5540" />
                    <RANKING order="4" place="4" resultid="5539" />
                    <RANKING order="5" place="5" resultid="5713" />
                    <RANKING order="6" place="6" resultid="5542" />
                    <RANKING order="7" place="7" resultid="5543" />
                    <RANKING order="8" place="8" resultid="5714" />
                    <RANKING order="9" place="9" resultid="5715" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4490" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5547" />
                    <RANKING order="2" place="2" resultid="5550" />
                    <RANKING order="3" place="3" resultid="5548" />
                    <RANKING order="4" place="4" resultid="5549" />
                    <RANKING order="5" place="5" resultid="5716" />
                    <RANKING order="6" place="6" resultid="5552" />
                    <RANKING order="7" place="7" resultid="5720" />
                    <RANKING order="8" place="8" resultid="5718" />
                    <RANKING order="9" place="9" resultid="5717" />
                    <RANKING order="10" place="10" resultid="5719" />
                    <RANKING order="11" place="-1" resultid="5551" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4491" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5721" />
                    <RANKING order="2" place="2" resultid="5722" />
                    <RANKING order="3" place="3" resultid="5557" />
                    <RANKING order="4" place="4" resultid="5559" />
                    <RANKING order="5" place="5" resultid="5560" />
                    <RANKING order="6" place="6" resultid="5558" />
                    <RANKING order="7" place="7" resultid="5726" />
                    <RANKING order="8" place="8" resultid="5724" />
                    <RANKING order="9" place="9" resultid="5723" />
                    <RANKING order="10" place="10" resultid="5562" />
                    <RANKING order="11" place="11" resultid="5561" />
                    <RANKING order="12" place="12" resultid="5727" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4792" agegroupid="4486" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4793" agegroupid="4486" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4794" agegroupid="4487" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4795" agegroupid="4487" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4796" agegroupid="4488" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4797" agegroupid="4488" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4798" agegroupid="4489" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4799" agegroupid="4489" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4800" agegroupid="4490" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4801" agegroupid="4490" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4802" agegroupid="4491" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4803" agegroupid="4491" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="4421" gender="M" number="6" order="15" round="FIN" preveventid="1089">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4462" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5463" />
                    <RANKING order="2" place="2" resultid="5464" />
                    <RANKING order="3" place="3" resultid="5465" />
                    <RANKING order="4" place="4" resultid="5466" />
                    <RANKING order="5" place="5" resultid="5467" />
                    <RANKING order="6" place="6" resultid="9024" />
                    <RANKING order="7" place="7" resultid="5468" />
                    <RANKING order="8" place="8" resultid="9022" />
                    <RANKING order="9" place="9" resultid="9023" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4463" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="9025" />
                    <RANKING order="2" place="2" resultid="5469" />
                    <RANKING order="3" place="3" resultid="5470" />
                    <RANKING order="4" place="4" resultid="5471" />
                    <RANKING order="5" place="5" resultid="5472" />
                    <RANKING order="6" place="6" resultid="5473" />
                    <RANKING order="7" place="7" resultid="5474" />
                    <RANKING order="8" place="8" resultid="9026" />
                    <RANKING order="9" place="9" resultid="9027" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4760" agegroupid="4462" final="F1" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9005" agegroupid="4462" final="F2" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4761" agegroupid="4463" final="F1" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9006" agegroupid="4463" final="F2" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="4425" gender="M" number="7" order="16" round="FIN" preveventid="4423">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4534" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5476" />
                    <RANKING order="2" place="2" resultid="5478" />
                    <RANKING order="3" place="3" resultid="5728" />
                    <RANKING order="4" place="4" resultid="5730" />
                    <RANKING order="5" place="5" resultid="5729" />
                    <RANKING order="6" place="-1" resultid="5479" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4535" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5603" />
                    <RANKING order="2" place="2" resultid="5731" />
                    <RANKING order="3" place="3" resultid="5732" />
                    <RANKING order="4" place="4" resultid="9034" />
                    <RANKING order="5" place="5" resultid="5605" />
                    <RANKING order="6" place="6" resultid="5604" />
                    <RANKING order="7" place="7" resultid="5733" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4536" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5736" />
                    <RANKING order="2" place="2" resultid="5734" />
                    <RANKING order="3" place="3" resultid="5535" />
                    <RANKING order="4" place="4" resultid="5537" />
                    <RANKING order="5" place="5" resultid="5536" />
                    <RANKING order="6" place="6" resultid="5735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4537" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5544" />
                    <RANKING order="2" place="2" resultid="5737" />
                    <RANKING order="3" place="3" resultid="10325" />
                    <RANKING order="4" place="4" resultid="5546" />
                    <RANKING order="5" place="5" resultid="5738" />
                    <RANKING order="6" place="6" resultid="5739" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4538" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5740" />
                    <RANKING order="2" place="2" resultid="5553" />
                    <RANKING order="3" place="3" resultid="5554" />
                    <RANKING order="4" place="4" resultid="5555" />
                    <RANKING order="5" place="5" resultid="5741" />
                    <RANKING order="6" place="6" resultid="5742" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4539" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5743" />
                    <RANKING order="2" place="2" resultid="5744" />
                    <RANKING order="3" place="3" resultid="5563" />
                    <RANKING order="4" place="4" resultid="5565" />
                    <RANKING order="5" place="5" resultid="5745" />
                    <RANKING order="6" place="6" resultid="10318" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4804" agegroupid="4534" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4805" agegroupid="4535" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4806" agegroupid="4536" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4807" agegroupid="4537" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4808" agegroupid="4538" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4809" agegroupid="4539" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="9999" agegroupid="4535" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1102" gender="M" number="8" order="17" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5271" agemax="9" agemin="9" name="[Colombo] Mirim 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2769" />
                    <RANKING order="2" place="2" resultid="3013" />
                    <RANKING order="3" place="3" resultid="1912" />
                    <RANKING order="4" place="4" resultid="4025" />
                    <RANKING order="5" place="5" resultid="2832" />
                    <RANKING order="6" place="6" resultid="2748" />
                    <RANKING order="7" place="7" resultid="3482" />
                    <RANKING order="8" place="8" resultid="2818" />
                    <RANKING order="9" place="9" resultid="2888" />
                    <RANKING order="10" place="10" resultid="3318" />
                    <RANKING order="11" place="11" resultid="2951" />
                    <RANKING order="12" place="12" resultid="2923" />
                    <RANKING order="13" place="13" resultid="2958" />
                    <RANKING order="14" place="14" resultid="2930" />
                    <RANKING order="15" place="-1" resultid="4227" />
                    <RANKING order="16" place="-1" resultid="2895" />
                    <RANKING order="17" place="-1" resultid="2909" />
                    <RANKING order="18" place="-1" resultid="2972" />
                    <RANKING order="19" place="-1" resultid="2985" />
                    <RANKING order="20" place="-1" resultid="2992" />
                    <RANKING order="21" place="-1" resultid="3061" />
                    <RANKING order="22" place="-1" resultid="3067" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5272" agemax="10" agemin="10" name="[Colombo] Mirim 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3425" />
                    <RANKING order="2" place="2" resultid="2692" />
                    <RANKING order="3" place="3" resultid="2881" />
                    <RANKING order="4" place="4" resultid="2589" />
                    <RANKING order="5" place="5" resultid="2596" />
                    <RANKING order="6" place="6" resultid="2657" />
                    <RANKING order="7" place="7" resultid="3963" />
                    <RANKING order="8" place="8" resultid="3020" />
                    <RANKING order="9" place="9" resultid="2582" />
                    <RANKING order="10" place="10" resultid="4073" />
                    <RANKING order="11" place="11" resultid="3970" />
                    <RANKING order="12" place="12" resultid="2685" />
                    <RANKING order="13" place="13" resultid="4101" />
                    <RANKING order="14" place="14" resultid="4094" />
                    <RANKING order="15" place="15" resultid="3990" />
                    <RANKING order="16" place="16" resultid="3074" />
                    <RANKING order="17" place="17" resultid="4122" />
                    <RANKING order="18" place="18" resultid="2664" />
                    <RANKING order="19" place="-1" resultid="1873" />
                    <RANKING order="20" place="-1" resultid="2624" />
                    <RANKING order="21" place="-1" resultid="2631" />
                    <RANKING order="22" place="-1" resultid="2650" />
                    <RANKING order="23" place="-1" resultid="2783" />
                    <RANKING order="24" place="-1" resultid="2804" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5273" agemax="9" agemin="9" name="[Maringá] Mirim 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3269" />
                    <RANKING order="2" place="2" resultid="1698" />
                    <RANKING order="3" place="3" resultid="1670" />
                    <RANKING order="4" place="4" resultid="1628" />
                    <RANKING order="5" place="5" resultid="1788" />
                    <RANKING order="6" place="6" resultid="3290" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5274" agemax="10" agemin="10" name="[Maringá] Mirim 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1621" />
                    <RANKING order="2" place="2" resultid="1684" />
                    <RANKING order="3" place="3" resultid="3432" />
                    <RANKING order="4" place="4" resultid="1710" />
                    <RANKING order="5" place="5" resultid="3343" />
                    <RANKING order="6" place="6" resultid="1745" />
                    <RANKING order="7" place="7" resultid="3398" />
                    <RANKING order="8" place="8" resultid="1663" />
                    <RANKING order="9" place="9" resultid="3439" />
                    <RANKING order="10" place="-1" resultid="1781" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4810" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4811" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4812" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4813" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4814" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4815" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4816" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4817" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4818" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4819" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4820" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1105" gender="M" number="9" order="18" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5313" agemax="11" agemin="11" name="[Colombo] Petiz 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1379" />
                    <RANKING order="2" place="2" resultid="2526" />
                    <RANKING order="3" place="3" resultid="2727" />
                    <RANKING order="4" place="4" resultid="3997" />
                    <RANKING order="5" place="5" resultid="3035" />
                    <RANKING order="6" place="6" resultid="4018" />
                    <RANKING order="7" place="7" resultid="2540" />
                    <RANKING order="8" place="8" resultid="2519" />
                    <RANKING order="9" place="9" resultid="2055" />
                    <RANKING order="10" place="10" resultid="3983" />
                    <RANKING order="11" place="11" resultid="2428" />
                    <RANKING order="12" place="12" resultid="3384" />
                    <RANKING order="13" place="13" resultid="2491" />
                    <RANKING order="14" place="14" resultid="2533" />
                    <RANKING order="15" place="15" resultid="4011" />
                    <RANKING order="16" place="16" resultid="2477" />
                    <RANKING order="17" place="17" resultid="4127" />
                    <RANKING order="18" place="18" resultid="3711" />
                    <RANKING order="19" place="19" resultid="3466" />
                    <RANKING order="20" place="20" resultid="3323" />
                    <RANKING order="21" place="-1" resultid="3049" />
                    <RANKING order="22" place="-1" resultid="3056" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5314" agemax="12" agemin="12" name="[Colombo] Petiz 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2311" />
                    <RANKING order="2" place="2" resultid="3677" />
                    <RANKING order="3" place="3" resultid="2358" />
                    <RANKING order="4" place="4" resultid="2346" />
                    <RANKING order="5" place="5" resultid="2365" />
                    <RANKING order="6" place="6" resultid="2339" />
                    <RANKING order="7" place="7" resultid="1866" />
                    <RANKING order="8" place="8" resultid="2393" />
                    <RANKING order="9" place="9" resultid="1919" />
                    <RANKING order="10" place="10" resultid="2318" />
                    <RANKING order="11" place="11" resultid="2414" />
                    <RANKING order="12" place="12" resultid="3942" />
                    <RANKING order="13" place="13" resultid="2400" />
                    <RANKING order="14" place="14" resultid="1834" />
                    <RANKING order="15" place="15" resultid="4087" />
                    <RANKING order="16" place="16" resultid="3905" />
                    <RANKING order="17" place="17" resultid="2554" />
                    <RANKING order="18" place="18" resultid="1828" />
                    <RANKING order="19" place="19" resultid="4148" />
                    <RANKING order="20" place="20" resultid="5260" />
                    <RANKING order="21" place="21" resultid="2353" />
                    <RANKING order="22" place="22" resultid="4046" />
                    <RANKING order="23" place="23" resultid="2505" />
                    <RANKING order="24" place="-1" resultid="4233" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5315" agemax="13" agemin="13" name="[Colombo] Infantil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2421" />
                    <RANKING order="2" place="2" resultid="1859" />
                    <RANKING order="3" place="3" resultid="3869" />
                    <RANKING order="4" place="4" resultid="4115" />
                    <RANKING order="5" place="5" resultid="3370" />
                    <RANKING order="6" place="6" resultid="2297" />
                    <RANKING order="7" place="7" resultid="2234" />
                    <RANKING order="8" place="8" resultid="2162" />
                    <RANKING order="9" place="9" resultid="3883" />
                    <RANKING order="10" place="10" resultid="3912" />
                    <RANKING order="11" place="11" resultid="2248" />
                    <RANKING order="12" place="12" resultid="3767" />
                    <RANKING order="13" place="13" resultid="2241" />
                    <RANKING order="14" place="14" resultid="1886" />
                    <RANKING order="15" place="15" resultid="3890" />
                    <RANKING order="16" place="16" resultid="3915" />
                    <RANKING order="17" place="17" resultid="2290" />
                    <RANKING order="18" place="18" resultid="2169" />
                    <RANKING order="19" place="19" resultid="2060" />
                    <RANKING order="20" place="20" resultid="2262" />
                    <RANKING order="21" place="21" resultid="2025" />
                    <RANKING order="22" place="-1" resultid="2561" />
                    <RANKING order="23" place="-1" resultid="3453" />
                    <RANKING order="24" place="-1" resultid="4134" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5316" agemax="14" agemin="14" name="[Colombo] Infantil 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2610" />
                    <RANKING order="2" place="2" resultid="2185" />
                    <RANKING order="3" place="3" resultid="2213" />
                    <RANKING order="4" place="4" resultid="2206" />
                    <RANKING order="5" place="5" resultid="4080" />
                    <RANKING order="6" place="6" resultid="4246" />
                    <RANKING order="7" place="7" resultid="2107" />
                    <RANKING order="8" place="8" resultid="2073" />
                    <RANKING order="9" place="9" resultid="2101" />
                    <RANKING order="10" place="10" resultid="2227" />
                    <RANKING order="11" place="11" resultid="4216" />
                    <RANKING order="12" place="12" resultid="4032" />
                    <RANKING order="13" place="13" resultid="3774" />
                    <RANKING order="14" place="-1" resultid="2220" />
                    <RANKING order="15" place="-1" resultid="3876" />
                    <RANKING order="16" place="-1" resultid="3897" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5317" agemax="15" agemin="15" name="[Colombo] Juvenil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4039" />
                    <RANKING order="2" place="2" resultid="3630" />
                    <RANKING order="3" place="3" resultid="3828" />
                    <RANKING order="4" place="4" resultid="1344" />
                    <RANKING order="5" place="5" resultid="3623" />
                    <RANKING order="6" place="6" resultid="1365" />
                    <RANKING order="7" place="7" resultid="2031" />
                    <RANKING order="8" place="8" resultid="2018" />
                    <RANKING order="9" place="9" resultid="3855" />
                    <RANKING order="10" place="10" resultid="4175" />
                    <RANKING order="11" place="11" resultid="2177" />
                    <RANKING order="12" place="-1" resultid="3835" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5318" agemax="-1" agemin="16" name="[Colombo] Juvenil 2/Sênior">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3329" />
                    <RANKING order="2" place="2" resultid="3618" />
                    <RANKING order="3" place="3" resultid="3637" />
                    <RANKING order="4" place="4" resultid="3816" />
                    <RANKING order="5" place="5" resultid="2085" />
                    <RANKING order="6" place="6" resultid="3848" />
                    <RANKING order="7" place="7" resultid="2148" />
                    <RANKING order="8" place="8" resultid="3704" />
                    <RANKING order="9" place="9" resultid="2134" />
                    <RANKING order="10" place="10" resultid="2011" />
                    <RANKING order="11" place="11" resultid="3336" />
                    <RANKING order="12" place="12" resultid="3788" />
                    <RANKING order="13" place="13" resultid="3690" />
                    <RANKING order="14" place="14" resultid="3670" />
                    <RANKING order="15" place="15" resultid="3684" />
                    <RANKING order="16" place="16" resultid="4202" />
                    <RANKING order="17" place="17" resultid="3795" />
                    <RANKING order="18" place="18" resultid="3658" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5319" agemax="11" agemin="11" name="[Maringá] Petiz 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1581" />
                    <RANKING order="2" place="2" resultid="1656" />
                    <RANKING order="3" place="3" resultid="1649" />
                    <RANKING order="4" place="4" resultid="1642" />
                    <RANKING order="5" place="5" resultid="1691" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5320" agemax="12" agemin="12" name="[Maringá] Petiz 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1588" />
                    <RANKING order="2" place="2" resultid="3136" />
                    <RANKING order="3" place="3" resultid="3562" />
                    <RANKING order="4" place="4" resultid="1574" />
                    <RANKING order="5" place="5" resultid="1595" />
                    <RANKING order="6" place="6" resultid="1553" />
                    <RANKING order="7" place="7" resultid="3220" />
                    <RANKING order="8" place="8" resultid="1635" />
                    <RANKING order="9" place="9" resultid="1427" />
                    <RANKING order="10" place="10" resultid="3503" />
                    <RANKING order="11" place="11" resultid="3582" />
                    <RANKING order="12" place="12" resultid="3595" />
                    <RANKING order="13" place="13" resultid="3589" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5321" agemax="13" agemin="13" name="[Maringá] Infantil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3164" />
                    <RANKING order="2" place="2" resultid="1407" />
                    <RANKING order="3" place="3" resultid="3192" />
                    <RANKING order="4" place="4" resultid="3108" />
                    <RANKING order="5" place="5" resultid="3171" />
                    <RANKING order="6" place="6" resultid="1455" />
                    <RANKING order="7" place="7" resultid="1992" />
                    <RANKING order="8" place="8" resultid="1462" />
                    <RANKING order="9" place="9" resultid="1985" />
                    <RANKING order="10" place="10" resultid="3122" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5322" agemax="14" agemin="14" name="[Maringá] Infantil 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1469" />
                    <RANKING order="2" place="2" resultid="3094" />
                    <RANKING order="3" place="3" resultid="3575" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5323" agemax="15" agemin="15" name="[Maringá] Juvenil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1420" />
                    <RANKING order="2" place="2" resultid="3536" />
                    <RANKING order="3" place="3" resultid="3157" />
                    <RANKING order="4" place="4" resultid="1441" />
                    <RANKING order="5" place="5" resultid="3509" />
                    <RANKING order="6" place="-1" resultid="1539" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5324" agemax="-1" agemin="16" name="[Maringá] Juvenil 2/Sênior">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1940" />
                    <RANKING order="2" place="2" resultid="1927" />
                    <RANKING order="3" place="3" resultid="1532" />
                    <RANKING order="4" place="4" resultid="1434" />
                    <RANKING order="5" place="5" resultid="1504" />
                    <RANKING order="6" place="6" resultid="1414" />
                    <RANKING order="7" place="7" resultid="1967" />
                    <RANKING order="8" place="8" resultid="3199" />
                    <RANKING order="9" place="9" resultid="3529" />
                    <RANKING order="10" place="10" resultid="1758" />
                    <RANKING order="11" place="11" resultid="1448" />
                    <RANKING order="12" place="12" resultid="3543" />
                    <RANKING order="13" place="13" resultid="3185" />
                    <RANKING order="14" place="14" resultid="1752" />
                    <RANKING order="15" place="-1" resultid="1476" />
                    <RANKING order="16" place="-1" resultid="1979" />
                    <RANKING order="17" place="-1" resultid="3515" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5253" order="1" status="OFFICIAL" />
                <HEAT heatid="4823" number="1" order="2" status="OFFICIAL" />
                <HEAT heatid="4824" number="2" order="3" status="OFFICIAL" />
                <HEAT heatid="4825" number="3" order="4" status="OFFICIAL" />
                <HEAT heatid="4826" number="4" order="5" status="OFFICIAL" />
                <HEAT heatid="4827" number="5" order="6" status="OFFICIAL" />
                <HEAT heatid="4828" number="6" order="7" status="OFFICIAL" />
                <HEAT heatid="4829" number="7" order="8" status="OFFICIAL" />
                <HEAT heatid="4830" number="8" order="9" status="OFFICIAL" />
                <HEAT heatid="4831" number="9" order="10" status="OFFICIAL" />
                <HEAT heatid="4832" number="10" order="11" status="OFFICIAL" />
                <HEAT heatid="4833" number="11" order="12" status="OFFICIAL" />
                <HEAT heatid="4834" number="12" order="13" status="OFFICIAL" />
                <HEAT heatid="4835" number="13" order="14" status="OFFICIAL" />
                <HEAT heatid="4836" number="14" order="15" status="OFFICIAL" />
                <HEAT heatid="4837" number="15" order="16" status="OFFICIAL" />
                <HEAT heatid="4838" number="16" order="17" status="OFFICIAL" />
                <HEAT heatid="4839" number="17" order="18" status="OFFICIAL" />
                <HEAT heatid="4840" number="18" order="19" status="OFFICIAL" />
                <HEAT heatid="4841" number="19" order="20" status="OFFICIAL" />
                <HEAT heatid="4842" number="20" order="21" status="OFFICIAL" />
                <HEAT heatid="4843" number="21" order="22" status="OFFICIAL" />
                <HEAT heatid="4844" number="22" order="23" status="OFFICIAL" />
                <HEAT heatid="4845" number="23" order="24" status="OFFICIAL" />
                <HEAT heatid="4846" number="24" order="25" status="OFFICIAL" />
                <HEAT heatid="4847" number="25" order="26" status="OFFICIAL" />
                <HEAT heatid="4848" number="26" order="27" status="OFFICIAL" />
                <HEAT heatid="4849" number="27" order="28" status="OFFICIAL" />
                <HEAT heatid="4850" number="28" order="29" status="OFFICIAL" />
                <HEAT heatid="4851" number="29" order="30" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="4429" gender="M" number="9" order="19" round="SEM" preveventid="1105">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4492" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5513" />
                    <RANKING order="2" place="2" resultid="5512" />
                    <RANKING order="3" place="3" resultid="5516" />
                    <RANKING order="4" place="4" resultid="5511" />
                    <RANKING order="5" place="5" resultid="5515" />
                    <RANKING order="6" place="6" resultid="5514" />
                    <RANKING order="7" place="7" resultid="5746" />
                    <RANKING order="8" place="8" resultid="5749" />
                    <RANKING order="9" place="9" resultid="5747" />
                    <RANKING order="10" place="10" resultid="5748" />
                    <RANKING order="11" place="11" resultid="5750" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4493" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5520" />
                    <RANKING order="2" place="2" resultid="5751" />
                    <RANKING order="3" place="3" resultid="5522" />
                    <RANKING order="4" place="4" resultid="5523" />
                    <RANKING order="5" place="5" resultid="5524" />
                    <RANKING order="6" place="6" resultid="5752" />
                    <RANKING order="7" place="7" resultid="5525" />
                    <RANKING order="8" place="8" resultid="5753" />
                    <RANKING order="9" place="9" resultid="5754" />
                    <RANKING order="10" place="10" resultid="5755" />
                    <RANKING order="11" place="11" resultid="5756" />
                    <RANKING order="12" place="-1" resultid="5521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4494" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5566" />
                    <RANKING order="2" place="2" resultid="5567" />
                    <RANKING order="3" place="3" resultid="5568" />
                    <RANKING order="4" place="4" resultid="5569" />
                    <RANKING order="5" place="5" resultid="5757" />
                    <RANKING order="6" place="6" resultid="5758" />
                    <RANKING order="7" place="7" resultid="5570" />
                    <RANKING order="8" place="8" resultid="5760" />
                    <RANKING order="9" place="9" resultid="5759" />
                    <RANKING order="10" place="10" resultid="5575" />
                    <RANKING order="11" place="11" resultid="5761" />
                    <RANKING order="12" place="12" resultid="5762" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4495" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5576" />
                    <RANKING order="2" place="2" resultid="5577" />
                    <RANKING order="3" place="3" resultid="5578" />
                    <RANKING order="4" place="4" resultid="5579" />
                    <RANKING order="5" place="5" resultid="5580" />
                    <RANKING order="6" place="6" resultid="5581" />
                    <RANKING order="7" place="7" resultid="5763" />
                    <RANKING order="8" place="8" resultid="5764" />
                    <RANKING order="9" place="9" resultid="5765" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4496" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5585" />
                    <RANKING order="2" place="2" resultid="5586" />
                    <RANKING order="3" place="3" resultid="5587" />
                    <RANKING order="4" place="4" resultid="5588" />
                    <RANKING order="5" place="5" resultid="5590" />
                    <RANKING order="6" place="6" resultid="5589" />
                    <RANKING order="7" place="7" resultid="5766" />
                    <RANKING order="8" place="8" resultid="5768" />
                    <RANKING order="9" place="9" resultid="5767" />
                    <RANKING order="10" place="10" resultid="5769" />
                    <RANKING order="11" place="11" resultid="5770" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4497" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5771" />
                    <RANKING order="2" place="2" resultid="5772" />
                    <RANKING order="3" place="3" resultid="5591" />
                    <RANKING order="4" place="4" resultid="5773" />
                    <RANKING order="5" place="5" resultid="5774" />
                    <RANKING order="6" place="6" resultid="5592" />
                    <RANKING order="7" place="7" resultid="5593" />
                    <RANKING order="8" place="8" resultid="5776" />
                    <RANKING order="9" place="9" resultid="5594" />
                    <RANKING order="10" place="10" resultid="5775" />
                    <RANKING order="11" place="11" resultid="5595" />
                    <RANKING order="12" place="12" resultid="5596" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4852" agegroupid="4492" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4853" agegroupid="4492" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4854" agegroupid="4493" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4855" agegroupid="4493" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4856" agegroupid="4494" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4857" agegroupid="4494" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4858" agegroupid="4495" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4859" agegroupid="4495" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4860" agegroupid="4496" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4861" agegroupid="4496" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4862" agegroupid="4497" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4863" agegroupid="4497" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="4427" gender="M" number="8" order="20" round="FIN" preveventid="1102">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4464" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5499" />
                    <RANKING order="2" place="2" resultid="5501" />
                    <RANKING order="3" place="3" resultid="5500" />
                    <RANKING order="4" place="4" resultid="5502" />
                    <RANKING order="5" place="5" resultid="9028" />
                    <RANKING order="6" place="6" resultid="9029" />
                    <RANKING order="7" place="7" resultid="10326" />
                    <RANKING order="8" place="8" resultid="9030" />
                    <RANKING order="9" place="9" resultid="5504" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4465" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5506" />
                    <RANKING order="2" place="2" resultid="5505" />
                    <RANKING order="3" place="3" resultid="5507" />
                    <RANKING order="4" place="4" resultid="9031" />
                    <RANKING order="5" place="5" resultid="5508" />
                    <RANKING order="6" place="6" resultid="5509" />
                    <RANKING order="7" place="7" resultid="9032" />
                    <RANKING order="8" place="8" resultid="5510" />
                    <RANKING order="9" place="9" resultid="9033" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4821" agegroupid="4464" final="F1" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="9007" agegroupid="4464" final="F2" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4822" agegroupid="4465" final="F1" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="9008" agegroupid="4465" final="F2" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="4431" gender="M" number="9" order="21" round="FIN" preveventid="4429">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4540" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5518" />
                    <RANKING order="2" place="2" resultid="5519" />
                    <RANKING order="3" place="3" resultid="5777" />
                    <RANKING order="4" place="4" resultid="5779" />
                    <RANKING order="5" place="5" resultid="5517" />
                    <RANKING order="6" place="6" resultid="5778" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4541" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5526" />
                    <RANKING order="2" place="2" resultid="5780" />
                    <RANKING order="3" place="3" resultid="5528" />
                    <RANKING order="4" place="4" resultid="5781" />
                    <RANKING order="5" place="5" resultid="5782" />
                    <RANKING order="6" place="6" resultid="5527" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4542" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5784" />
                    <RANKING order="2" place="2" resultid="5783" />
                    <RANKING order="3" place="3" resultid="5572" />
                    <RANKING order="4" place="4" resultid="5574" />
                    <RANKING order="5" place="5" resultid="5573" />
                    <RANKING order="6" place="6" resultid="5785" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4543" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5582" />
                    <RANKING order="2" place="2" resultid="5786" />
                    <RANKING order="3" place="3" resultid="5584" />
                    <RANKING order="4" place="4" resultid="5583" />
                    <RANKING order="5" place="5" resultid="5787" />
                    <RANKING order="6" place="6" resultid="5788" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4544" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5600" />
                    <RANKING order="2" place="2" resultid="5789" />
                    <RANKING order="3" place="3" resultid="5601" />
                    <RANKING order="4" place="4" resultid="5790" />
                    <RANKING order="5" place="5" resultid="5602" />
                    <RANKING order="6" place="6" resultid="5791" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4545" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5792" />
                    <RANKING order="2" place="2" resultid="5793" />
                    <RANKING order="3" place="3" resultid="5794" />
                    <RANKING order="4" place="4" resultid="5597" />
                    <RANKING order="5" place="5" resultid="5599" />
                    <RANKING order="6" place="6" resultid="5598" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4864" agegroupid="4540" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4865" agegroupid="4541" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4866" agegroupid="4542" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4867" agegroupid="4543" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4868" agegroupid="4544" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4869" agegroupid="4545" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1115" gender="M" number="10" order="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="8" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1116" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4259" />
                    <RANKING order="2" place="2" resultid="1803" />
                    <RANKING order="3" place="3" resultid="3085" />
                    <RANKING order="4" place="4" resultid="3494" />
                    <RANKING order="5" place="5" resultid="3606" />
                    <RANKING order="6" place="-1" resultid="3081" />
                    <RANKING order="7" place="-1" resultid="2121" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4870" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4871" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5251" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-12-07" daytime="15:10" endtime="03:44" number="2" officialmeeting="14:30" warmupfrom="14:30" warmupuntil="15:00">
          <EVENTS>
            <EVENT eventid="1117" gender="F" number="11" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4605" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1769" />
                    <RANKING order="2" place="2" resultid="3026" />
                    <RANKING order="3" place="3" resultid="2091" />
                    <RANKING order="4" place="4" resultid="1798" />
                    <RANKING order="5" place="5" resultid="3030" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4872" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4873" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1119" gender="F" number="12" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5916" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2436" />
                    <RANKING order="2" place="2" resultid="2485" />
                    <RANKING order="3" place="3" resultid="3249" />
                    <RANKING order="4" place="4" resultid="2499" />
                    <RANKING order="5" place="-1" resultid="1547" />
                    <RANKING order="6" place="-1" resultid="3242" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5917" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2513" />
                    <RANKING order="2" place="2" resultid="2457" />
                    <RANKING order="3" place="3" resultid="1561" />
                    <RANKING order="4" place="4" resultid="3950" />
                    <RANKING order="5" place="5" resultid="4109" />
                    <RANKING order="6" place="6" resultid="3923" />
                    <RANKING order="7" place="7" resultid="3235" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5918" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2305" />
                    <RANKING order="2" place="2" resultid="2284" />
                    <RANKING order="3" place="3" resultid="2277" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5919" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1814" />
                    <RANKING order="2" place="2" resultid="2193" />
                    <RANKING order="3" place="3" resultid="1961" />
                    <RANKING order="4" place="4" resultid="4196" />
                    <RANKING order="5" place="-1" resultid="3719" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5920" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1519" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5921" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3652" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4874" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4875" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4876" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4877" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4878" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1129" gender="F" number="13" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5959" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2826" />
                    <RANKING order="2" place="2" resultid="2791" />
                    <RANKING order="3" place="3" resultid="2812" />
                    <RANKING order="4" place="4" resultid="1394" />
                    <RANKING order="5" place="5" resultid="1775" />
                    <RANKING order="6" place="6" resultid="2763" />
                    <RANKING order="7" place="7" resultid="2756" />
                    <RANKING order="8" place="8" resultid="3298" />
                    <RANKING order="9" place="9" resultid="2777" />
                    <RANKING order="10" place="-1" resultid="2854" />
                    <RANKING order="11" place="-1" resultid="2917" />
                    <RANKING order="12" place="-1" resultid="2938" />
                    <RANKING order="13" place="-1" resultid="2980" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5958" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3930" />
                    <RANKING order="2" place="2" resultid="2569" />
                    <RANKING order="3" place="3" resultid="2735" />
                    <RANKING order="4" place="4" resultid="4169" />
                    <RANKING order="5" place="5" resultid="4067" />
                    <RANKING order="6" place="6" resultid="2721" />
                    <RANKING order="7" place="7" resultid="4210" />
                    <RANKING order="8" place="8" resultid="2576" />
                    <RANKING order="9" place="9" resultid="2742" />
                    <RANKING order="10" place="10" resultid="1615" />
                    <RANKING order="11" place="11" resultid="3256" />
                    <RANKING order="12" place="12" resultid="1718" />
                    <RANKING order="13" place="13" resultid="3392" />
                    <RANKING order="14" place="14" resultid="2679" />
                    <RANKING order="15" place="15" resultid="3602" />
                    <RANKING order="16" place="-1" resultid="4155" />
                    <RANKING order="17" place="-1" resultid="2639" />
                    <RANKING order="18" place="-1" resultid="2700" />
                    <RANKING order="19" place="-1" resultid="3000" />
                    <RANKING order="20" place="-1" resultid="3474" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5952" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2443" />
                    <RANKING order="2" place="2" resultid="3312" />
                    <RANKING order="3" place="3" resultid="2966" />
                    <RANKING order="4" place="4" resultid="2548" />
                    <RANKING order="5" place="5" resultid="1568" />
                    <RANKING order="6" place="6" resultid="2714" />
                    <RANKING order="7" place="7" resultid="4054" />
                    <RANKING order="8" place="-1" resultid="3488" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5953" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2373" />
                    <RANKING order="2" place="2" resultid="3116" />
                    <RANKING order="3" place="3" resultid="2408" />
                    <RANKING order="4" place="4" resultid="1601" />
                    <RANKING order="5" place="5" resultid="2387" />
                    <RANKING order="6" place="6" resultid="3207" />
                    <RANKING order="7" place="7" resultid="2380" />
                    <RANKING order="8" place="8" resultid="1880" />
                    <RANKING order="9" place="9" resultid="4142" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5954" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2256" />
                    <RANKING order="2" place="2" resultid="2875" />
                    <RANKING order="3" place="3" resultid="2270" />
                    <RANKING order="4" place="4" resultid="3151" />
                    <RANKING order="5" place="5" resultid="3284" />
                    <RANKING order="6" place="6" resultid="1974" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5955" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3612" />
                    <RANKING order="2" place="2" resultid="2604" />
                    <RANKING order="3" place="3" resultid="2200" />
                    <RANKING order="4" place="4" resultid="3409" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5956" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2038" />
                    <RANKING order="2" place="2" resultid="1359" />
                    <RANKING order="3" place="3" resultid="3102" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5957" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1512" />
                    <RANKING order="2" place="2" resultid="3740" />
                    <RANKING order="3" place="3" resultid="3822" />
                    <RANKING order="4" place="4" resultid="3523" />
                    <RANKING order="5" place="-1" resultid="1822" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4879" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4880" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4881" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4882" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4883" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4884" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4885" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4886" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4887" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4888" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4889" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4890" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1141" gender="F" number="14" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5911" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2092" />
                    <RANKING order="2" place="2" resultid="3027" />
                    <RANKING order="3" place="3" resultid="1770" />
                    <RANKING order="4" place="4" resultid="3031" />
                    <RANKING order="5" place="5" resultid="1799" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4891" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4892" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1143" gender="F" number="15" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5922" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3278" />
                    <RANKING order="2" place="2" resultid="4240" />
                    <RANKING order="3" place="3" resultid="3378" />
                    <RANKING order="4" place="4" resultid="1853" />
                    <RANKING order="5" place="5" resultid="2618" />
                    <RANKING order="6" place="6" resultid="1608" />
                    <RANKING order="7" place="7" resultid="3699" />
                    <RANKING order="8" place="8" resultid="1569" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5923" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2334" />
                    <RANKING order="2" place="2" resultid="2327" />
                    <RANKING order="3" place="3" resultid="2471" />
                    <RANKING order="4" place="4" resultid="2945" />
                    <RANKING order="5" place="5" resultid="2708" />
                    <RANKING order="6" place="6" resultid="3951" />
                    <RANKING order="7" place="7" resultid="3783" />
                    <RANKING order="8" place="8" resultid="3549" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5924" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2868" />
                    <RANKING order="2" place="2" resultid="1491" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5925" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1484" />
                    <RANKING order="2" place="2" resultid="3645" />
                    <RANKING order="3" place="3" resultid="1809" />
                    <RANKING order="4" place="4" resultid="3180" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5926" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2143" />
                    <RANKING order="2" place="2" resultid="1954" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5927" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1947" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4893" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4894" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4895" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4896" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4897" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1153" gender="F" number="16" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5960" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2827" />
                    <RANKING order="2" place="2" resultid="2792" />
                    <RANKING order="3" place="3" resultid="2841" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5961" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2570" />
                    <RANKING order="2" place="2" resultid="4061" />
                    <RANKING order="3" place="3" resultid="3228" />
                    <RANKING order="4" place="4" resultid="2673" />
                    <RANKING order="5" place="5" resultid="4156" />
                    <RANKING order="6" place="-1" resultid="2861" />
                    <RANKING order="7" place="-1" resultid="1719" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5962" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3957" />
                    <RANKING order="2" place="2" resultid="3250" />
                    <RANKING order="3" place="3" resultid="3277" />
                    <RANKING order="4" place="4" resultid="3263" />
                    <RANKING order="5" place="5" resultid="3214" />
                    <RANKING order="6" place="6" resultid="4005" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5963" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2514" />
                    <RANKING order="2" place="2" resultid="3145" />
                    <RANKING order="3" place="3" resultid="2388" />
                    <RANKING order="4" place="4" resultid="3352" />
                    <RANKING order="5" place="5" resultid="2080" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5964" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2285" />
                    <RANKING order="2" place="2" resultid="1498" />
                    <RANKING order="3" place="3" resultid="2278" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5965" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1934" />
                    <RANKING order="2" place="2" resultid="2194" />
                    <RANKING order="3" place="3" resultid="3727" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5966" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3805" />
                    <RANKING order="2" place="-1" resultid="1526" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5967" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3733" />
                    <RANKING order="2" place="2" resultid="3359" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4898" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4899" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4900" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4901" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4902" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4903" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1165" gender="F" number="17" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5968" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3747" />
                    <RANKING order="2" place="2" resultid="2847" />
                    <RANKING order="3" place="3" resultid="3754" />
                    <RANKING order="4" place="4" resultid="3043" />
                    <RANKING order="5" place="5" resultid="1894" />
                    <RANKING order="6" place="6" resultid="2764" />
                    <RANKING order="7" place="7" resultid="2813" />
                    <RANKING order="8" place="8" resultid="2840" />
                    <RANKING order="9" place="9" resultid="2778" />
                    <RANKING order="10" place="-1" resultid="2757" />
                    <RANKING order="11" place="-1" resultid="2855" />
                    <RANKING order="12" place="-1" resultid="2903" />
                    <RANKING order="13" place="-1" resultid="2918" />
                    <RANKING order="14" place="-1" resultid="2939" />
                    <RANKING order="15" place="-1" resultid="3007" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5969" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4060" />
                    <RANKING order="2" place="2" resultid="1725" />
                    <RANKING order="3" place="3" resultid="4170" />
                    <RANKING order="4" place="4" resultid="2672" />
                    <RANKING order="5" place="5" resultid="2577" />
                    <RANKING order="6" place="6" resultid="4068" />
                    <RANKING order="7" place="7" resultid="2798" />
                    <RANKING order="8" place="8" resultid="4211" />
                    <RANKING order="9" place="9" resultid="2736" />
                    <RANKING order="10" place="10" resultid="2722" />
                    <RANKING order="11" place="11" resultid="2743" />
                    <RANKING order="12" place="12" resultid="3556" />
                    <RANKING order="13" place="13" resultid="3257" />
                    <RANKING order="14" place="14" resultid="2680" />
                    <RANKING order="15" place="15" resultid="3761" />
                    <RANKING order="16" place="16" resultid="3447" />
                    <RANKING order="17" place="-1" resultid="2701" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5970" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2437" />
                    <RANKING order="2" place="2" resultid="2486" />
                    <RANKING order="3" place="3" resultid="2500" />
                    <RANKING order="4" place="4" resultid="3243" />
                    <RANKING order="5" place="5" resultid="2049" />
                    <RANKING order="6" place="6" resultid="3698" />
                    <RANKING order="7" place="7" resultid="3130" />
                    <RANKING order="8" place="8" resultid="4183" />
                    <RANKING order="9" place="-1" resultid="3489" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5971" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2333" />
                    <RANKING order="2" place="2" resultid="2326" />
                    <RANKING order="3" place="3" resultid="2707" />
                    <RANKING order="4" place="4" resultid="2458" />
                    <RANKING order="5" place="5" resultid="1562" />
                    <RANKING order="6" place="6" resultid="2079" />
                    <RANKING order="7" place="7" resultid="3782" />
                    <RANKING order="8" place="8" resultid="1373" />
                    <RANKING order="9" place="9" resultid="3416" />
                    <RANKING order="10" place="10" resultid="3305" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5972" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2450" />
                    <RANKING order="2" place="2" resultid="1387" />
                    <RANKING order="3" place="3" resultid="3152" />
                    <RANKING order="4" place="4" resultid="3285" />
                    <RANKING order="5" place="5" resultid="4162" />
                    <RANKING order="6" place="-1" resultid="1901" />
                    <RANKING order="7" place="-1" resultid="2156" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5973" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1815" />
                    <RANKING order="2" place="2" resultid="1962" />
                    <RANKING order="3" place="3" resultid="4197" />
                    <RANKING order="4" place="4" resultid="4189" />
                    <RANKING order="5" place="5" resultid="3179" />
                    <RANKING order="6" place="6" resultid="3720" />
                    <RANKING order="7" place="7" resultid="3726" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5974" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1352" />
                    <RANKING order="2" place="2" resultid="3804" />
                    <RANKING order="3" place="3" resultid="3103" />
                    <RANKING order="4" place="4" resultid="3863" />
                    <RANKING order="5" place="-1" resultid="1520" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5975" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3653" />
                    <RANKING order="2" place="2" resultid="1841" />
                    <RANKING order="3" place="3" resultid="3664" />
                    <RANKING order="4" place="4" resultid="2067" />
                    <RANKING order="5" place="5" resultid="4254" />
                    <RANKING order="6" place="-1" resultid="1765" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4904" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4905" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4906" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4907" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4908" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4909" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4910" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4911" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4912" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4913" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4914" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4915" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="4916" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="4917" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1177" gender="F" number="18" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5912" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3028" />
                    <RANKING order="2" place="2" resultid="2093" />
                    <RANKING order="3" place="3" resultid="1771" />
                    <RANKING order="4" place="4" resultid="1800" />
                    <RANKING order="5" place="5" resultid="3032" />
                    <RANKING order="6" place="6" resultid="3479" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4918" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4919" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1179" gender="F" number="19" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5928" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1678" />
                    <RANKING order="2" place="2" resultid="2444" />
                    <RANKING order="3" place="3" resultid="3313" />
                    <RANKING order="4" place="4" resultid="2464" />
                    <RANKING order="5" place="5" resultid="2967" />
                    <RANKING order="6" place="6" resultid="2549" />
                    <RANKING order="7" place="7" resultid="2715" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5929" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2374" />
                    <RANKING order="2" place="2" resultid="3117" />
                    <RANKING order="3" place="3" resultid="2409" />
                    <RANKING order="4" place="4" resultid="3144" />
                    <RANKING order="5" place="5" resultid="1602" />
                    <RANKING order="6" place="6" resultid="3351" />
                    <RANKING order="7" place="7" resultid="1881" />
                    <RANKING order="8" place="-1" resultid="4110" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5930" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2257" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5931" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3613" />
                    <RANKING order="2" place="2" resultid="3410" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5932" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1360" />
                    <RANKING order="2" place="2" resultid="2142" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5933" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3823" />
                    <RANKING order="2" place="2" resultid="3358" />
                    <RANKING order="3" place="3" resultid="3524" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4920" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4921" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4922" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4923" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1189" gender="F" number="20" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5976" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3748" />
                    <RANKING order="2" place="2" resultid="2848" />
                    <RANKING order="3" place="3" resultid="3755" />
                    <RANKING order="4" place="4" resultid="3044" />
                    <RANKING order="5" place="5" resultid="1776" />
                    <RANKING order="6" place="6" resultid="1895" />
                    <RANKING order="7" place="7" resultid="3299" />
                    <RANKING order="8" place="-1" resultid="2904" />
                    <RANKING order="9" place="-1" resultid="2981" />
                    <RANKING order="10" place="-1" resultid="3008" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5977" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3931" />
                    <RANKING order="2" place="2" resultid="3229" />
                    <RANKING order="3" place="3" resultid="2862" />
                    <RANKING order="4" place="4" resultid="1726" />
                    <RANKING order="5" place="5" resultid="2799" />
                    <RANKING order="6" place="6" resultid="1616" />
                    <RANKING order="7" place="7" resultid="3448" />
                    <RANKING order="8" place="8" resultid="2000" />
                    <RANKING order="9" place="9" resultid="3557" />
                    <RANKING order="10" place="10" resultid="3762" />
                    <RANKING order="11" place="11" resultid="3393" />
                    <RANKING order="12" place="12" resultid="3603" />
                    <RANKING order="13" place="-1" resultid="1731" />
                    <RANKING order="14" place="-1" resultid="2640" />
                    <RANKING order="15" place="-1" resultid="3001" />
                    <RANKING order="16" place="-1" resultid="3475" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5978" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3958" />
                    <RANKING order="2" place="2" resultid="1679" />
                    <RANKING order="3" place="3" resultid="2465" />
                    <RANKING order="4" place="4" resultid="4241" />
                    <RANKING order="5" place="5" resultid="1854" />
                    <RANKING order="6" place="6" resultid="3379" />
                    <RANKING order="7" place="7" resultid="2050" />
                    <RANKING order="8" place="8" resultid="4006" />
                    <RANKING order="9" place="9" resultid="3264" />
                    <RANKING order="10" place="10" resultid="2619" />
                    <RANKING order="11" place="11" resultid="3215" />
                    <RANKING order="12" place="12" resultid="3131" />
                    <RANKING order="13" place="13" resultid="1609" />
                    <RANKING order="14" place="14" resultid="3365" />
                    <RANKING order="15" place="-1" resultid="1548" />
                    <RANKING order="16" place="-1" resultid="3937" />
                    <RANKING order="17" place="-1" resultid="3978" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5979" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2472" />
                    <RANKING order="2" place="2" resultid="2381" />
                    <RANKING order="3" place="3" resultid="2946" />
                    <RANKING order="4" place="4" resultid="3461" />
                    <RANKING order="5" place="5" resultid="3924" />
                    <RANKING order="6" place="6" resultid="3208" />
                    <RANKING order="7" place="7" resultid="1374" />
                    <RANKING order="8" place="8" resultid="3550" />
                    <RANKING order="9" place="9" resultid="3417" />
                    <RANKING order="10" place="10" resultid="3236" />
                    <RANKING order="11" place="11" resultid="4143" />
                    <RANKING order="12" place="12" resultid="3306" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5980" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2451" />
                    <RANKING order="2" place="2" resultid="1388" />
                    <RANKING order="3" place="3" resultid="2876" />
                    <RANKING order="4" place="4" resultid="2869" />
                    <RANKING order="5" place="5" resultid="1492" />
                    <RANKING order="6" place="6" resultid="2306" />
                    <RANKING order="7" place="7" resultid="2271" />
                    <RANKING order="8" place="8" resultid="4163" />
                    <RANKING order="9" place="9" resultid="1499" />
                    <RANKING order="10" place="10" resultid="1902" />
                    <RANKING order="11" place="-1" resultid="2157" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5981" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1816" />
                    <RANKING order="2" place="2" resultid="1485" />
                    <RANKING order="3" place="3" resultid="2201" />
                    <RANKING order="4" place="4" resultid="2605" />
                    <RANKING order="5" place="5" resultid="3646" />
                    <RANKING order="6" place="6" resultid="1935" />
                    <RANKING order="7" place="7" resultid="4190" />
                    <RANKING order="8" place="8" resultid="1810" />
                    <RANKING order="9" place="9" resultid="3570" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5982" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3806" />
                    <RANKING order="2" place="2" resultid="3843" />
                    <RANKING order="3" place="3" resultid="1353" />
                    <RANKING order="4" place="4" resultid="1955" />
                    <RANKING order="5" place="5" resultid="3864" />
                    <RANKING order="6" place="-1" resultid="1527" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5983" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3741" />
                    <RANKING order="2" place="2" resultid="1823" />
                    <RANKING order="3" place="3" resultid="1513" />
                    <RANKING order="4" place="4" resultid="1948" />
                    <RANKING order="5" place="5" resultid="3734" />
                    <RANKING order="6" place="6" resultid="3665" />
                    <RANKING order="7" place="7" resultid="1842" />
                    <RANKING order="8" place="8" resultid="2068" />
                    <RANKING order="9" place="9" resultid="1766" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4924" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4925" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4926" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4927" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4928" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4929" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4930" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4931" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4932" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4933" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4934" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4935" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="4936" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="4937" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="4938" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="4939" number="16" order="16" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1201" gender="M" number="21" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5913" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1794" />
                    <RANKING order="2" place="2" resultid="2112" />
                    <RANKING order="3" place="3" resultid="1740" />
                    <RANKING order="4" place="4" resultid="3404" />
                    <RANKING order="5" place="5" resultid="4222" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4940" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4941" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1203" gender="M" number="22" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5934" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2527" />
                    <RANKING order="2" place="2" resultid="3984" />
                    <RANKING order="3" place="3" resultid="1657" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5935" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2312" />
                    <RANKING order="2" place="2" resultid="3678" />
                    <RANKING order="3" place="3" resultid="1589" />
                    <RANKING order="4" place="4" resultid="2366" />
                    <RANKING order="5" place="5" resultid="2340" />
                    <RANKING order="6" place="6" resultid="3137" />
                    <RANKING order="7" place="7" resultid="3221" />
                    <RANKING order="8" place="8" resultid="2415" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5936" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3165" />
                    <RANKING order="2" place="2" resultid="3870" />
                    <RANKING order="3" place="3" resultid="3371" />
                    <RANKING order="4" place="4" resultid="1463" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5937" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1470" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5938" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1345" />
                    <RANKING order="2" place="2" resultid="3624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5939" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1533" />
                    <RANKING order="2" place="2" resultid="3330" />
                    <RANKING order="3" place="3" resultid="3530" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4942" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4943" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4944" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4945" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1213" gender="M" number="23" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5984" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2749" />
                    <RANKING order="2" place="2" resultid="2931" />
                    <RANKING order="3" place="3" resultid="1699" />
                    <RANKING order="4" place="4" resultid="4026" />
                    <RANKING order="5" place="5" resultid="1629" />
                    <RANKING order="6" place="6" resultid="1671" />
                    <RANKING order="7" place="7" resultid="2819" />
                    <RANKING order="8" place="8" resultid="2952" />
                    <RANKING order="9" place="9" resultid="2959" />
                    <RANKING order="10" place="-1" resultid="2896" />
                    <RANKING order="11" place="-1" resultid="2986" />
                    <RANKING order="12" place="-1" resultid="3062" />
                    <RANKING order="13" place="-1" resultid="3068" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5985" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1622" />
                    <RANKING order="2" place="2" resultid="2597" />
                    <RANKING order="3" place="3" resultid="2693" />
                    <RANKING order="4" place="4" resultid="3971" />
                    <RANKING order="5" place="5" resultid="2686" />
                    <RANKING order="6" place="6" resultid="2583" />
                    <RANKING order="7" place="7" resultid="3344" />
                    <RANKING order="8" place="8" resultid="3433" />
                    <RANKING order="9" place="9" resultid="4074" />
                    <RANKING order="10" place="10" resultid="3021" />
                    <RANKING order="11" place="11" resultid="4095" />
                    <RANKING order="12" place="12" resultid="4102" />
                    <RANKING order="13" place="13" resultid="2658" />
                    <RANKING order="14" place="14" resultid="3399" />
                    <RANKING order="15" place="15" resultid="1664" />
                    <RANKING order="16" place="16" resultid="3440" />
                    <RANKING order="17" place="17" resultid="3075" />
                    <RANKING order="18" place="-1" resultid="1782" />
                    <RANKING order="19" place="-1" resultid="2632" />
                    <RANKING order="20" place="-1" resultid="2651" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5986" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3036" />
                    <RANKING order="2" place="2" resultid="3998" />
                    <RANKING order="3" place="3" resultid="1643" />
                    <RANKING order="4" place="4" resultid="2534" />
                    <RANKING order="5" place="5" resultid="3050" />
                    <RANKING order="6" place="-1" resultid="4128" />
                    <RANKING order="7" place="-1" resultid="2478" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5987" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2359" />
                    <RANKING order="2" place="2" resultid="2394" />
                    <RANKING order="3" place="3" resultid="2555" />
                    <RANKING order="4" place="4" resultid="1554" />
                    <RANKING order="5" place="5" resultid="1428" />
                    <RANKING order="6" place="6" resultid="1835" />
                    <RANKING order="7" place="7" resultid="3583" />
                    <RANKING order="8" place="8" resultid="3590" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5988" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2249" />
                    <RANKING order="2" place="2" resultid="2291" />
                    <RANKING order="3" place="3" resultid="1456" />
                    <RANKING order="4" place="4" resultid="3884" />
                    <RANKING order="5" place="5" resultid="2263" />
                    <RANKING order="6" place="-1" resultid="2242" />
                    <RANKING order="7" place="-1" resultid="3123" />
                    <RANKING order="8" place="-1" resultid="3454" />
                    <RANKING order="9" place="-1" resultid="4135" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5989" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3095" />
                    <RANKING order="2" place="2" resultid="2102" />
                    <RANKING order="3" place="3" resultid="4247" />
                    <RANKING order="4" place="4" resultid="2214" />
                    <RANKING order="5" place="5" resultid="2207" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5990" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3856" />
                    <RANKING order="2" place="2" resultid="2019" />
                    <RANKING order="3" place="3" resultid="1442" />
                    <RANKING order="4" place="4" resultid="3537" />
                    <RANKING order="5" place="-1" resultid="2032" />
                    <RANKING order="6" place="-1" resultid="3631" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5991" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1415" />
                    <RANKING order="2" place="2" resultid="1534" />
                    <RANKING order="3" place="3" resultid="1980" />
                    <RANKING order="4" place="4" resultid="3789" />
                    <RANKING order="5" place="5" resultid="3685" />
                    <RANKING order="6" place="6" resultid="3705" />
                    <RANKING order="7" place="7" resultid="1759" />
                    <RANKING order="8" place="8" resultid="3186" />
                    <RANKING order="9" place="-1" resultid="3516" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4946" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4947" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4948" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4949" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4950" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4951" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4952" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4953" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4954" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4955" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4956" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4957" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="4958" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="4959" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1225" gender="M" number="24" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5914" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1795" />
                    <RANKING order="2" place="2" resultid="2113" />
                    <RANKING order="3" place="3" resultid="1741" />
                    <RANKING order="4" place="4" resultid="4223" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4960" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4961" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1227" gender="M" number="25" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5940" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2541" />
                    <RANKING order="2" place="2" resultid="3385" />
                    <RANKING order="3" place="3" resultid="1582" />
                    <RANKING order="4" place="4" resultid="2492" />
                    <RANKING order="5" place="5" resultid="1650" />
                    <RANKING order="6" place="6" resultid="3712" />
                    <RANKING order="7" place="7" resultid="3467" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5941" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2313" />
                    <RANKING order="2" place="2" resultid="2347" />
                    <RANKING order="3" place="3" resultid="3679" />
                    <RANKING order="4" place="4" resultid="1829" />
                    <RANKING order="5" place="5" resultid="1636" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5942" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2422" />
                    <RANKING order="2" place="2" resultid="1408" />
                    <RANKING order="3" place="3" resultid="2163" />
                    <RANKING order="4" place="4" resultid="2235" />
                    <RANKING order="5" place="5" resultid="3768" />
                    <RANKING order="6" place="6" resultid="3916" />
                    <RANKING order="7" place="7" resultid="3891" />
                    <RANKING order="8" place="8" resultid="1993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5943" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2186" />
                    <RANKING order="2" place="2" resultid="2611" />
                    <RANKING order="3" place="3" resultid="4217" />
                    <RANKING order="4" place="4" resultid="2221" />
                    <RANKING order="5" place="5" resultid="4033" />
                    <RANKING order="6" place="6" resultid="3576" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5944" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1346" />
                    <RANKING order="2" place="2" resultid="3158" />
                    <RANKING order="3" place="3" resultid="4176" />
                    <RANKING order="4" place="4" resultid="2178" />
                    <RANKING order="5" place="-1" resultid="3836" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5945" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3638" />
                    <RANKING order="2" place="2" resultid="2012" />
                    <RANKING order="3" place="3" resultid="3849" />
                    <RANKING order="4" place="4" resultid="1435" />
                    <RANKING order="5" place="5" resultid="3817" />
                    <RANKING order="6" place="6" resultid="2086" />
                    <RANKING order="7" place="7" resultid="3796" />
                    <RANKING order="8" place="8" resultid="4203" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4962" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4963" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4964" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4965" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4966" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4967" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4968" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5254" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1237" gender="M" number="26" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5992" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2771" />
                    <RANKING order="2" place="2" resultid="3291" />
                    <RANKING order="3" place="3" resultid="1700" />
                    <RANKING order="4" place="4" resultid="2820" />
                    <RANKING order="5" place="5" resultid="1789" />
                    <RANKING order="6" place="6" resultid="2890" />
                    <RANKING order="7" place="-1" resultid="2834" />
                    <RANKING order="8" place="-1" resultid="2932" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5993" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2591" />
                    <RANKING order="2" place="2" resultid="2687" />
                    <RANKING order="3" place="3" resultid="2883" />
                    <RANKING order="4" place="-1" resultid="2806" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5994" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1380" />
                    <RANKING order="2" place="2" resultid="2429" />
                    <RANKING order="3" place="3" resultid="2520" />
                    <RANKING order="4" place="4" resultid="4019" />
                    <RANKING order="5" place="5" resultid="1658" />
                    <RANKING order="6" place="6" resultid="2479" />
                    <RANKING order="7" place="7" resultid="1651" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5995" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1575" />
                    <RANKING order="2" place="2" resultid="1590" />
                    <RANKING order="3" place="3" resultid="2401" />
                    <RANKING order="4" place="4" resultid="2319" />
                    <RANKING order="5" place="5" resultid="4047" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5996" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4116" />
                    <RANKING order="2" place="2" resultid="3871" />
                    <RANKING order="3" place="3" resultid="3166" />
                    <RANKING order="4" place="4" resultid="3172" />
                    <RANKING order="5" place="5" resultid="2243" />
                    <RANKING order="6" place="6" resultid="2299" />
                    <RANKING order="7" place="7" resultid="2170" />
                    <RANKING order="8" place="8" resultid="1986" />
                    <RANKING order="9" place="9" resultid="3110" />
                    <RANKING order="10" place="-1" resultid="2562" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5997" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3877" />
                    <RANKING order="2" place="2" resultid="2228" />
                    <RANKING order="3" place="3" resultid="4034" />
                    <RANKING order="4" place="4" resultid="3775" />
                    <RANKING order="5" place="5" resultid="2215" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5998" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1421" />
                    <RANKING order="2" place="2" resultid="3830" />
                    <RANKING order="3" place="3" resultid="1366" />
                    <RANKING order="4" place="4" resultid="3625" />
                    <RANKING order="5" place="-1" resultid="1540" />
                    <RANKING order="6" place="-1" resultid="4041" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5999" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3691" />
                    <RANKING order="2" place="2" resultid="1505" />
                    <RANKING order="3" place="3" resultid="3200" />
                    <RANKING order="4" place="4" resultid="3671" />
                    <RANKING order="5" place="5" resultid="3337" />
                    <RANKING order="6" place="6" resultid="2149" />
                    <RANKING order="7" place="-1" resultid="1941" />
                    <RANKING order="8" place="-1" resultid="1477" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4969" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4970" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4971" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4972" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4973" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4974" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4975" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4976" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4977" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1249" gender="M" number="27" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6000" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1913" />
                    <RANKING order="2" place="2" resultid="2770" />
                    <RANKING order="3" place="3" resultid="3270" />
                    <RANKING order="4" place="4" resultid="2750" />
                    <RANKING order="5" place="5" resultid="2924" />
                    <RANKING order="6" place="6" resultid="2889" />
                    <RANKING order="7" place="7" resultid="2953" />
                    <RANKING order="8" place="8" resultid="2960" />
                    <RANKING order="9" place="-1" resultid="2833" />
                    <RANKING order="10" place="-1" resultid="2897" />
                    <RANKING order="11" place="-1" resultid="2910" />
                    <RANKING order="12" place="-1" resultid="2973" />
                    <RANKING order="13" place="-1" resultid="2993" />
                    <RANKING order="14" place="-1" resultid="3014" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6001" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2882" />
                    <RANKING order="2" place="2" resultid="2694" />
                    <RANKING order="3" place="3" resultid="3426" />
                    <RANKING order="4" place="4" resultid="2590" />
                    <RANKING order="5" place="5" resultid="2598" />
                    <RANKING order="6" place="6" resultid="1685" />
                    <RANKING order="7" place="7" resultid="3964" />
                    <RANKING order="8" place="8" resultid="3434" />
                    <RANKING order="9" place="9" resultid="4075" />
                    <RANKING order="10" place="10" resultid="2659" />
                    <RANKING order="11" place="11" resultid="2584" />
                    <RANKING order="12" place="12" resultid="1711" />
                    <RANKING order="13" place="13" resultid="3022" />
                    <RANKING order="14" place="14" resultid="1746" />
                    <RANKING order="15" place="15" resultid="3991" />
                    <RANKING order="16" place="16" resultid="2665" />
                    <RANKING order="17" place="-1" resultid="1783" />
                    <RANKING order="18" place="-1" resultid="2625" />
                    <RANKING order="19" place="-1" resultid="2652" />
                    <RANKING order="20" place="-1" resultid="2784" />
                    <RANKING order="21" place="-1" resultid="2805" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6002" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2528" />
                    <RANKING order="2" place="2" resultid="2728" />
                    <RANKING order="3" place="3" resultid="1583" />
                    <RANKING order="4" place="4" resultid="3985" />
                    <RANKING order="5" place="5" resultid="3386" />
                    <RANKING order="6" place="6" resultid="3713" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6003" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1867" />
                    <RANKING order="2" place="2" resultid="2360" />
                    <RANKING order="3" place="3" resultid="3138" />
                    <RANKING order="4" place="4" resultid="2341" />
                    <RANKING order="5" place="5" resultid="3563" />
                    <RANKING order="6" place="6" resultid="1920" />
                    <RANKING order="7" place="7" resultid="3943" />
                    <RANKING order="8" place="8" resultid="1836" />
                    <RANKING order="9" place="9" resultid="4088" />
                    <RANKING order="10" place="10" resultid="2506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6004" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1860" />
                    <RANKING order="2" place="2" resultid="3193" />
                    <RANKING order="3" place="3" resultid="3372" />
                    <RANKING order="4" place="4" resultid="2298" />
                    <RANKING order="5" place="5" resultid="3109" />
                    <RANKING order="6" place="6" resultid="1887" />
                    <RANKING order="7" place="7" resultid="2264" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6005" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1471" />
                    <RANKING order="2" place="2" resultid="2208" />
                    <RANKING order="3" place="3" resultid="4081" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6006" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4040" />
                    <RANKING order="2" place="2" resultid="3632" />
                    <RANKING order="3" place="3" resultid="3829" />
                    <RANKING order="4" place="4" resultid="3159" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6007" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1928" />
                    <RANKING order="2" place="2" resultid="3331" />
                    <RANKING order="3" place="3" resultid="2135" />
                    <RANKING order="4" place="4" resultid="3531" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4978" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4979" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4980" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4981" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4982" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4983" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4984" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4985" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4986" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4987" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4988" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4989" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1261" gender="M" number="28" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5915" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1796" />
                    <RANKING order="2" place="2" resultid="1742" />
                    <RANKING order="3" place="3" resultid="2114" />
                    <RANKING order="4" place="4" resultid="3405" />
                    <RANKING order="5" place="5" resultid="4224" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4990" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4991" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1263" gender="M" number="29" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5946" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3037" />
                    <RANKING order="2" place="2" resultid="3999" />
                    <RANKING order="3" place="3" resultid="1644" />
                    <RANKING order="4" place="4" resultid="4012" />
                    <RANKING order="5" place="5" resultid="2535" />
                    <RANKING order="6" place="6" resultid="1692" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5947" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2395" />
                    <RANKING order="2" place="2" resultid="3906" />
                    <RANKING order="3" place="3" resultid="2556" />
                    <RANKING order="4" place="4" resultid="1429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5948" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2292" />
                    <RANKING order="2" place="2" resultid="3769" />
                    <RANKING order="3" place="3" resultid="3885" />
                    <RANKING order="4" place="4" resultid="3173" />
                    <RANKING order="5" place="5" resultid="1457" />
                    <RANKING order="6" place="-1" resultid="3455" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5949" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3096" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5950" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5951" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1449" />
                    <RANKING order="2" place="2" resultid="3201" />
                    <RANKING order="3" place="3" resultid="3187" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4992" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4993" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4994" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4995" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1273" gender="M" number="30" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6008" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4027" />
                    <RANKING order="2" place="2" resultid="1914" />
                    <RANKING order="3" place="3" resultid="3015" />
                    <RANKING order="4" place="4" resultid="3271" />
                    <RANKING order="5" place="5" resultid="1790" />
                    <RANKING order="6" place="6" resultid="1672" />
                    <RANKING order="7" place="7" resultid="1630" />
                    <RANKING order="8" place="8" resultid="3292" />
                    <RANKING order="9" place="9" resultid="4228" />
                    <RANKING order="10" place="-1" resultid="2911" />
                    <RANKING order="11" place="-1" resultid="2925" />
                    <RANKING order="12" place="-1" resultid="2974" />
                    <RANKING order="13" place="-1" resultid="2987" />
                    <RANKING order="14" place="-1" resultid="2994" />
                    <RANKING order="15" place="-1" resultid="3063" />
                    <RANKING order="16" place="-1" resultid="3069" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6009" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1623" />
                    <RANKING order="2" place="2" resultid="3427" />
                    <RANKING order="3" place="3" resultid="1686" />
                    <RANKING order="4" place="4" resultid="3972" />
                    <RANKING order="5" place="5" resultid="3345" />
                    <RANKING order="6" place="6" resultid="3992" />
                    <RANKING order="7" place="7" resultid="1712" />
                    <RANKING order="8" place="8" resultid="3965" />
                    <RANKING order="9" place="9" resultid="4103" />
                    <RANKING order="10" place="10" resultid="4096" />
                    <RANKING order="11" place="11" resultid="1747" />
                    <RANKING order="12" place="12" resultid="3400" />
                    <RANKING order="13" place="13" resultid="1665" />
                    <RANKING order="14" place="14" resultid="3076" />
                    <RANKING order="15" place="15" resultid="2666" />
                    <RANKING order="16" place="16" resultid="3441" />
                    <RANKING order="17" place="-1" resultid="1874" />
                    <RANKING order="18" place="-1" resultid="2626" />
                    <RANKING order="19" place="-1" resultid="2633" />
                    <RANKING order="20" place="-1" resultid="2785" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6010" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1381" />
                    <RANKING order="2" place="2" resultid="2729" />
                    <RANKING order="3" place="3" resultid="4020" />
                    <RANKING order="4" place="4" resultid="2521" />
                    <RANKING order="5" place="5" resultid="2542" />
                    <RANKING order="6" place="6" resultid="2430" />
                    <RANKING order="7" place="7" resultid="4013" />
                    <RANKING order="8" place="8" resultid="2493" />
                    <RANKING order="9" place="9" resultid="1693" />
                    <RANKING order="10" place="10" resultid="3468" />
                    <RANKING order="11" place="11" resultid="3324" />
                    <RANKING order="12" place="12" resultid="3051" />
                    <RANKING order="13" place="-1" resultid="4129" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6011" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1576" />
                    <RANKING order="2" place="2" resultid="3907" />
                    <RANKING order="3" place="3" resultid="2348" />
                    <RANKING order="4" place="4" resultid="1868" />
                    <RANKING order="5" place="5" resultid="2367" />
                    <RANKING order="6" place="6" resultid="2320" />
                    <RANKING order="7" place="7" resultid="1555" />
                    <RANKING order="8" place="8" resultid="3222" />
                    <RANKING order="9" place="9" resultid="2416" />
                    <RANKING order="10" place="10" resultid="2402" />
                    <RANKING order="11" place="11" resultid="1830" />
                    <RANKING order="12" place="12" resultid="3944" />
                    <RANKING order="13" place="13" resultid="3564" />
                    <RANKING order="14" place="14" resultid="1921" />
                    <RANKING order="15" place="15" resultid="1637" />
                    <RANKING order="16" place="16" resultid="4048" />
                    <RANKING order="17" place="17" resultid="4089" />
                    <RANKING order="18" place="18" resultid="3584" />
                    <RANKING order="19" place="19" resultid="4149" />
                    <RANKING order="20" place="20" resultid="3504" />
                    <RANKING order="21" place="21" resultid="2507" />
                    <RANKING order="22" place="22" resultid="3596" />
                    <RANKING order="23" place="-1" resultid="4234" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6012" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1409" />
                    <RANKING order="2" place="2" resultid="2423" />
                    <RANKING order="3" place="3" resultid="1861" />
                    <RANKING order="4" place="4" resultid="2250" />
                    <RANKING order="5" place="5" resultid="4117" />
                    <RANKING order="6" place="6" resultid="2164" />
                    <RANKING order="7" place="7" resultid="2236" />
                    <RANKING order="8" place="8" resultid="3917" />
                    <RANKING order="9" place="9" resultid="2061" />
                    <RANKING order="10" place="10" resultid="3194" />
                    <RANKING order="11" place="11" resultid="3892" />
                    <RANKING order="12" place="12" resultid="1888" />
                    <RANKING order="13" place="13" resultid="2171" />
                    <RANKING order="14" place="14" resultid="1987" />
                    <RANKING order="15" place="15" resultid="1994" />
                    <RANKING order="16" place="16" resultid="1464" />
                    <RANKING order="17" place="17" resultid="2026" />
                    <RANKING order="18" place="18" resultid="3124" />
                    <RANKING order="19" place="-1" resultid="2563" />
                    <RANKING order="20" place="-1" resultid="4136" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6013" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2612" />
                    <RANKING order="2" place="2" resultid="2187" />
                    <RANKING order="3" place="3" resultid="4218" />
                    <RANKING order="4" place="4" resultid="2229" />
                    <RANKING order="5" place="5" resultid="3878" />
                    <RANKING order="6" place="6" resultid="2222" />
                    <RANKING order="7" place="7" resultid="4248" />
                    <RANKING order="8" place="8" resultid="3776" />
                    <RANKING order="9" place="9" resultid="4082" />
                    <RANKING order="10" place="10" resultid="3577" />
                    <RANKING order="11" place="-1" resultid="2108" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6014" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1422" />
                    <RANKING order="2" place="2" resultid="3857" />
                    <RANKING order="3" place="3" resultid="4177" />
                    <RANKING order="4" place="4" resultid="1367" />
                    <RANKING order="5" place="5" resultid="2020" />
                    <RANKING order="6" place="6" resultid="3538" />
                    <RANKING order="7" place="7" resultid="3510" />
                    <RANKING order="8" place="8" resultid="2179" />
                    <RANKING order="9" place="-1" resultid="1541" />
                    <RANKING order="10" place="-1" resultid="3837" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6015" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1968" />
                    <RANKING order="2" place="2" resultid="3809" />
                    <RANKING order="3" place="3" resultid="3692" />
                    <RANKING order="4" place="4" resultid="3850" />
                    <RANKING order="5" place="5" resultid="3639" />
                    <RANKING order="6" place="6" resultid="2013" />
                    <RANKING order="7" place="7" resultid="1436" />
                    <RANKING order="8" place="8" resultid="3818" />
                    <RANKING order="9" place="9" resultid="3706" />
                    <RANKING order="10" place="10" resultid="3790" />
                    <RANKING order="11" place="11" resultid="1506" />
                    <RANKING order="12" place="12" resultid="2087" />
                    <RANKING order="13" place="13" resultid="3338" />
                    <RANKING order="14" place="14" resultid="2136" />
                    <RANKING order="15" place="15" resultid="3672" />
                    <RANKING order="16" place="16" resultid="1450" />
                    <RANKING order="17" place="17" resultid="2150" />
                    <RANKING order="18" place="18" resultid="1760" />
                    <RANKING order="19" place="19" resultid="3797" />
                    <RANKING order="20" place="20" resultid="4204" />
                    <RANKING order="21" place="21" resultid="1753" />
                    <RANKING order="22" place="-1" resultid="1478" />
                    <RANKING order="23" place="-1" resultid="3517" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4996" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4997" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4998" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4999" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5000" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5001" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5002" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5003" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5004" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="5005" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="5006" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="5007" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="5008" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="5009" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="5010" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="5011" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="5012" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="5013" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="5014" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="5015" number="20" order="20" status="OFFICIAL" />
                <HEAT heatid="5016" number="21" order="21" status="OFFICIAL" />
                <HEAT heatid="5017" number="22" order="22" status="OFFICIAL" />
                <HEAT heatid="5018" number="23" order="23" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-12-08" daytime="08:10" endtime="12:22" number="3" officialmeeting="07:30" warmupfrom="07:30" warmupuntil="08:00">
          <POOL lanemin="1" lanemax="8" />
          <EVENTS>
            <EVENT eventid="1298" gender="F" number="31" order="1" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5813" agemax="9" agemin="9" name="[Colombo] Mirim 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2828" />
                    <RANKING order="2" place="2" resultid="3749" />
                    <RANKING order="3" place="3" resultid="2793" />
                    <RANKING order="4" place="4" resultid="2814" />
                    <RANKING order="5" place="5" resultid="1395" />
                    <RANKING order="6" place="6" resultid="2849" />
                    <RANKING order="7" place="7" resultid="2765" />
                    <RANKING order="8" place="8" resultid="2758" />
                    <RANKING order="9" place="9" resultid="3756" />
                    <RANKING order="10" place="10" resultid="2842" />
                    <RANKING order="11" place="11" resultid="1896" />
                    <RANKING order="12" place="12" resultid="2779" />
                    <RANKING order="13" place="-1" resultid="2856" />
                    <RANKING order="14" place="-1" resultid="2905" />
                    <RANKING order="15" place="-1" resultid="2919" />
                    <RANKING order="16" place="-1" resultid="2940" />
                    <RANKING order="17" place="-1" resultid="2982" />
                    <RANKING order="18" place="-1" resultid="3009" />
                    <RANKING order="19" place="-1" resultid="3045" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5814" agemax="10" agemin="10" name="[Colombo] Mirim 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3932" />
                    <RANKING order="2" place="2" resultid="2571" />
                    <RANKING order="3" place="3" resultid="4062" />
                    <RANKING order="4" place="4" resultid="2863" />
                    <RANKING order="5" place="5" resultid="2737" />
                    <RANKING order="6" place="6" resultid="2744" />
                    <RANKING order="7" place="7" resultid="2723" />
                    <RANKING order="8" place="8" resultid="2674" />
                    <RANKING order="9" place="9" resultid="4069" />
                    <RANKING order="10" place="10" resultid="4157" />
                    <RANKING order="11" place="11" resultid="2578" />
                    <RANKING order="12" place="12" resultid="2097" />
                    <RANKING order="13" place="13" resultid="1400" />
                    <RANKING order="14" place="14" resultid="2800" />
                    <RANKING order="15" place="15" resultid="2681" />
                    <RANKING order="16" place="16" resultid="3763" />
                    <RANKING order="17" place="-1" resultid="2641" />
                    <RANKING order="18" place="-1" resultid="2702" />
                    <RANKING order="19" place="-1" resultid="3002" />
                    <RANKING order="20" place="-1" resultid="4171" />
                    <RANKING order="21" place="-1" resultid="4212" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5815" agemax="9" agemin="9" name="[Maringá] Mirim 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1777" />
                    <RANKING order="2" place="2" resultid="3300" />
                    <RANKING order="3" place="3" resultid="1737" />
                    <RANKING order="4" place="4" resultid="1706" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5816" agemax="10" agemin="10" name="[Maringá] Mirim 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3230" />
                    <RANKING order="2" place="2" resultid="1727" />
                    <RANKING order="3" place="3" resultid="1617" />
                    <RANKING order="4" place="4" resultid="3258" />
                    <RANKING order="5" place="5" resultid="3394" />
                    <RANKING order="6" place="6" resultid="2001" />
                    <RANKING order="7" place="7" resultid="1720" />
                    <RANKING order="8" place="8" resultid="3558" />
                    <RANKING order="9" place="9" resultid="3604" />
                    <RANKING order="10" place="10" resultid="3449" />
                    <RANKING order="11" place="-1" resultid="1732" />
                    <RANKING order="12" place="-1" resultid="3476" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5020" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5021" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5023" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5024" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5025" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5026" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5027" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="5028" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1301" gender="F" number="32" order="2" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5829" agemax="11" agemin="11" name="[Colombo] Petiz 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2551" />
                    <RANKING order="2" place="2" resultid="2969" />
                    <RANKING order="3" place="3" resultid="2467" />
                    <RANKING order="4" place="4" resultid="2446" />
                    <RANKING order="5" place="5" resultid="3381" />
                    <RANKING order="6" place="6" resultid="2621" />
                    <RANKING order="7" place="7" resultid="3280" />
                    <RANKING order="8" place="8" resultid="3960" />
                    <RANKING order="9" place="9" resultid="4243" />
                    <RANKING order="10" place="10" resultid="2488" />
                    <RANKING order="11" place="11" resultid="3939" />
                    <RANKING order="12" place="12" resultid="2717" />
                    <RANKING order="13" place="13" resultid="3980" />
                    <RANKING order="14" place="14" resultid="2502" />
                    <RANKING order="15" place="15" resultid="1909" />
                    <RANKING order="16" place="16" resultid="3701" />
                    <RANKING order="17" place="17" resultid="2052" />
                    <RANKING order="18" place="18" resultid="2647" />
                    <RANKING order="19" place="19" resultid="4008" />
                    <RANKING order="20" place="20" resultid="1856" />
                    <RANKING order="21" place="21" resultid="3367" />
                    <RANKING order="22" place="22" resultid="4185" />
                    <RANKING order="23" place="-1" resultid="4056" />
                    <RANKING order="24" place="-1" resultid="2439" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5830" agemax="12" agemin="12" name="[Colombo] Petiz 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2376" />
                    <RANKING order="2" place="2" resultid="4112" />
                    <RANKING order="3" place="3" resultid="2336" />
                    <RANKING order="4" place="4" resultid="2329" />
                    <RANKING order="5" place="5" resultid="2411" />
                    <RANKING order="6" place="6" resultid="2516" />
                    <RANKING order="7" place="7" resultid="2948" />
                    <RANKING order="8" place="8" resultid="2390" />
                    <RANKING order="9" place="9" resultid="3926" />
                    <RANKING order="10" place="10" resultid="2710" />
                    <RANKING order="11" place="11" resultid="2383" />
                    <RANKING order="12" place="12" resultid="2474" />
                    <RANKING order="13" place="13" resultid="2460" />
                    <RANKING order="14" place="14" resultid="3354" />
                    <RANKING order="15" place="15" resultid="3953" />
                    <RANKING order="16" place="16" resultid="1883" />
                    <RANKING order="17" place="17" resultid="3463" />
                    <RANKING order="18" place="18" resultid="1849" />
                    <RANKING order="19" place="19" resultid="3785" />
                    <RANKING order="20" place="20" resultid="2082" />
                    <RANKING order="21" place="21" resultid="4145" />
                    <RANKING order="22" place="22" resultid="1376" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5831" agemax="13" agemin="13" name="[Colombo] Infantil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2259" />
                    <RANKING order="2" place="2" resultid="2878" />
                    <RANKING order="3" place="3" resultid="2453" />
                    <RANKING order="4" place="4" resultid="2273" />
                    <RANKING order="5" place="5" resultid="2280" />
                    <RANKING order="6" place="6" resultid="2308" />
                    <RANKING order="7" place="7" resultid="3154" />
                    <RANKING order="8" place="8" resultid="2871" />
                    <RANKING order="9" place="9" resultid="2287" />
                    <RANKING order="10" place="10" resultid="2159" />
                    <RANKING order="11" place="11" resultid="1390" />
                    <RANKING order="12" place="12" resultid="1904" />
                    <RANKING order="13" place="13" resultid="4165" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5832" agemax="14" agemin="14" name="[Colombo] Infantil 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2607" />
                    <RANKING order="2" place="2" resultid="3615" />
                    <RANKING order="3" place="3" resultid="2196" />
                    <RANKING order="4" place="4" resultid="2203" />
                    <RANKING order="5" place="5" resultid="1818" />
                    <RANKING order="6" place="6" resultid="3412" />
                    <RANKING order="7" place="7" resultid="3648" />
                    <RANKING order="8" place="8" resultid="4199" />
                    <RANKING order="9" place="9" resultid="1812" />
                    <RANKING order="10" place="10" resultid="4192" />
                    <RANKING order="11" place="11" resultid="3729" />
                    <RANKING order="12" place="12" resultid="3722" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5833" agemax="15" agemin="15" name="[Colombo] Juvenil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2040" />
                    <RANKING order="2" place="2" resultid="1362" />
                    <RANKING order="3" place="3" resultid="1355" />
                    <RANKING order="4" place="4" resultid="2008" />
                    <RANKING order="5" place="5" resultid="2145" />
                    <RANKING order="6" place="6" resultid="2045" />
                    <RANKING order="7" place="7" resultid="3866" />
                    <RANKING order="8" place="-1" resultid="3845" />
                    <RANKING order="9" place="-1" resultid="3105" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5834" agemax="-1" agemin="16" name="[Colombo] Juvenil 2/Sênior">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1825" />
                    <RANKING order="2" place="2" resultid="3743" />
                    <RANKING order="3" place="3" resultid="3736" />
                    <RANKING order="4" place="4" resultid="3825" />
                    <RANKING order="5" place="5" resultid="3655" />
                    <RANKING order="6" place="6" resultid="4256" />
                    <RANKING order="7" place="7" resultid="3667" />
                    <RANKING order="8" place="8" resultid="2070" />
                    <RANKING order="9" place="-1" resultid="1844" />
                    <RANKING order="10" place="-1" resultid="3361" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5835" agemax="11" agemin="11" name="[Maringá] Petiz 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3315" />
                    <RANKING order="2" place="2" resultid="3252" />
                    <RANKING order="3" place="3" resultid="1571" />
                    <RANKING order="4" place="4" resultid="3217" />
                    <RANKING order="5" place="5" resultid="3133" />
                    <RANKING order="6" place="6" resultid="3245" />
                    <RANKING order="7" place="7" resultid="3266" />
                    <RANKING order="8" place="8" resultid="1611" />
                    <RANKING order="9" place="9" resultid="3491" />
                    <RANKING order="10" place="-1" resultid="1681" />
                    <RANKING order="11" place="-1" resultid="1550" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5836" agemax="12" agemin="12" name="[Maringá] Petiz 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3119" />
                    <RANKING order="2" place="2" resultid="3210" />
                    <RANKING order="3" place="3" resultid="3147" />
                    <RANKING order="4" place="4" resultid="1604" />
                    <RANKING order="5" place="5" resultid="1564" />
                    <RANKING order="6" place="6" resultid="3238" />
                    <RANKING order="7" place="7" resultid="3552" />
                    <RANKING order="8" place="8" resultid="3308" />
                    <RANKING order="9" place="-1" resultid="3419" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5837" agemax="13" agemin="13" name="[Maringá] Infantil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3287" />
                    <RANKING order="2" place="2" resultid="1494" />
                    <RANKING order="3" place="3" resultid="1976" />
                    <RANKING order="4" place="4" resultid="1501" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5838" agemax="14" agemin="14" name="[Maringá] Infantil 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3182" />
                    <RANKING order="2" place="2" resultid="1487" />
                    <RANKING order="3" place="3" resultid="1937" />
                    <RANKING order="4" place="4" resultid="1964" />
                    <RANKING order="5" place="5" resultid="3572" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5839" agemax="15" agemin="15" name="[Maringá] Juvenil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1957" />
                    <RANKING order="2" place="2" resultid="1522" />
                    <RANKING order="3" place="-1" resultid="1529" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5840" agemax="-1" agemin="16" name="[Maringá] Juvenil 2/Sênior">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1515" />
                    <RANKING order="2" place="2" resultid="3526" />
                    <RANKING order="3" place="3" resultid="1950" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5031" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5032" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5033" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5034" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5036" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5037" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5038" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5040" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5041" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="5042" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="5044" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="5045" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="5046" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="5047" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="5048" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="5049" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="5050" number="20" order="20" status="OFFICIAL" />
                <HEAT heatid="5051" number="21" order="21" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="4433" gender="F" number="31" order="3" round="FIN" preveventid="1298">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4466" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10080" />
                    <RANKING order="2" place="2" resultid="10081" />
                    <RANKING order="3" place="3" resultid="10082" />
                    <RANKING order="4" place="4" resultid="10083" />
                    <RANKING order="5" place="5" resultid="10084" />
                    <RANKING order="6" place="6" resultid="10078" />
                    <RANKING order="7" place="7" resultid="10001" />
                    <RANKING order="8" place="8" resultid="10002" />
                    <RANKING order="9" place="9" resultid="10004" />
                    <RANKING order="10" place="10" resultid="10003" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4467" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10085" />
                    <RANKING order="2" place="2" resultid="10087" />
                    <RANKING order="3" place="3" resultid="10086" />
                    <RANKING order="4" place="4" resultid="10090" />
                    <RANKING order="5" place="5" resultid="10005" />
                    <RANKING order="6" place="6" resultid="10088" />
                    <RANKING order="7" place="7" resultid="10089" />
                    <RANKING order="8" place="8" resultid="10006" />
                    <RANKING order="9" place="9" resultid="10008" />
                    <RANKING order="10" place="10" resultid="10007" />
                    <RANKING order="11" place="11" resultid="10009" />
                    <RANKING order="12" place="12" resultid="10010" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5029" agegroupid="4466" final="F1" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5030" agegroupid="4466" final="F2" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6064" agegroupid="4467" final="F1" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6065" agegroupid="4467" final="F2" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5801" gender="F" number="32" order="4" round="FIN" preveventid="1301">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5883" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10092" />
                    <RANKING order="2" place="2" resultid="10011" />
                    <RANKING order="3" place="3" resultid="10091" />
                    <RANKING order="4" place="4" resultid="10093" />
                    <RANKING order="5" place="5" resultid="10094" />
                    <RANKING order="6" place="6" resultid="10095" />
                    <RANKING order="7" place="7" resultid="10096" />
                    <RANKING order="8" place="8" resultid="10012" />
                    <RANKING order="9" place="9" resultid="10013" />
                    <RANKING order="10" place="10" resultid="10014" />
                    <RANKING order="11" place="11" resultid="10015" />
                    <RANKING order="12" place="12" resultid="10016" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5884" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10017" />
                    <RANKING order="2" place="2" resultid="10097" />
                    <RANKING order="3" place="3" resultid="10098" />
                    <RANKING order="4" place="4" resultid="10102" />
                    <RANKING order="5" place="5" resultid="10099" />
                    <RANKING order="6" place="6" resultid="10101" />
                    <RANKING order="7" place="7" resultid="10100" />
                    <RANKING order="8" place="8" resultid="10019" />
                    <RANKING order="9" place="9" resultid="10018" />
                    <RANKING order="10" place="10" resultid="10020" />
                    <RANKING order="11" place="11" resultid="10021" />
                    <RANKING order="12" place="12" resultid="10022" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5885" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10155" />
                    <RANKING order="2" place="2" resultid="10154" />
                    <RANKING order="3" place="3" resultid="10156" />
                    <RANKING order="4" place="4" resultid="10157" />
                    <RANKING order="5" place="5" resultid="10160" />
                    <RANKING order="6" place="6" resultid="10158" />
                    <RANKING order="7" place="7" resultid="10023" />
                    <RANKING order="8" place="8" resultid="10025" />
                    <RANKING order="9" place="9" resultid="10024" />
                    <RANKING order="10" place="-1" resultid="10026" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5886" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10104" />
                    <RANKING order="2" place="2" resultid="10103" />
                    <RANKING order="3" place="3" resultid="10108" />
                    <RANKING order="4" place="4" resultid="10105" />
                    <RANKING order="5" place="5" resultid="10106" />
                    <RANKING order="6" place="6" resultid="10107" />
                    <RANKING order="7" place="7" resultid="10027" />
                    <RANKING order="8" place="8" resultid="10028" />
                    <RANKING order="9" place="9" resultid="10029" />
                    <RANKING order="10" place="10" resultid="10030" />
                    <RANKING order="11" place="-1" resultid="10031" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5887" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10161" />
                    <RANKING order="2" place="2" resultid="10162" />
                    <RANKING order="3" place="3" resultid="10163" />
                    <RANKING order="4" place="4" resultid="10327" />
                    <RANKING order="5" place="5" resultid="10544" />
                    <RANKING order="6" place="6" resultid="10033" />
                    <RANKING order="7" place="7" resultid="10166" />
                    <RANKING order="8" place="8" resultid="10034" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5888" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10036" />
                    <RANKING order="2" place="2" resultid="10168" />
                    <RANKING order="3" place="3" resultid="10167" />
                    <RANKING order="4" place="4" resultid="10170" />
                    <RANKING order="5" place="5" resultid="10169" />
                    <RANKING order="6" place="6" resultid="10037" />
                    <RANKING order="7" place="7" resultid="10171" />
                    <RANKING order="8" place="8" resultid="10172" />
                    <RANKING order="9" place="9" resultid="10038" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6066" agegroupid="5883" final="F1" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6067" agegroupid="5883" final="F2" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6068" agegroupid="5884" final="F1" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6069" agegroupid="5884" final="F2" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6070" agegroupid="5885" final="F1" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6071" agegroupid="5885" final="F2" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6072" agegroupid="5886" final="F1" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6073" agegroupid="5886" final="F2" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6074" agegroupid="5887" final="F1" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6075" agegroupid="5887" final="F2" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6076" agegroupid="5888" final="F1" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="6077" agegroupid="5888" final="F2" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1311" gender="F" number="33" order="5" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5817" agemax="9" agemin="9" name="[Colombo] Mirim 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3750" />
                    <RANKING order="2" place="2" resultid="2850" />
                    <RANKING order="3" place="3" resultid="2794" />
                    <RANKING order="4" place="4" resultid="2829" />
                    <RANKING order="5" place="5" resultid="3757" />
                    <RANKING order="6" place="6" resultid="2766" />
                    <RANKING order="7" place="7" resultid="1396" />
                    <RANKING order="8" place="8" resultid="1897" />
                    <RANKING order="9" place="9" resultid="3046" />
                    <RANKING order="10" place="10" resultid="2815" />
                    <RANKING order="11" place="11" resultid="2843" />
                    <RANKING order="12" place="12" resultid="2759" />
                    <RANKING order="13" place="13" resultid="2780" />
                    <RANKING order="14" place="-1" resultid="2857" />
                    <RANKING order="15" place="-1" resultid="2906" />
                    <RANKING order="16" place="-1" resultid="2920" />
                    <RANKING order="17" place="-1" resultid="2941" />
                    <RANKING order="18" place="-1" resultid="2983" />
                    <RANKING order="19" place="-1" resultid="3010" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5818" agemax="10" agemin="10" name="[Colombo] Mirim 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4063" />
                    <RANKING order="2" place="2" resultid="3933" />
                    <RANKING order="3" place="3" resultid="2572" />
                    <RANKING order="4" place="4" resultid="2864" />
                    <RANKING order="5" place="5" resultid="2675" />
                    <RANKING order="6" place="6" resultid="1401" />
                    <RANKING order="7" place="7" resultid="2682" />
                    <RANKING order="8" place="8" resultid="2745" />
                    <RANKING order="9" place="9" resultid="4070" />
                    <RANKING order="10" place="10" resultid="2724" />
                    <RANKING order="11" place="11" resultid="2579" />
                    <RANKING order="12" place="12" resultid="4158" />
                    <RANKING order="13" place="13" resultid="2801" />
                    <RANKING order="14" place="14" resultid="2738" />
                    <RANKING order="15" place="15" resultid="3764" />
                    <RANKING order="16" place="16" resultid="2098" />
                    <RANKING order="17" place="-1" resultid="2642" />
                    <RANKING order="18" place="-1" resultid="2703" />
                    <RANKING order="19" place="-1" resultid="3003" />
                    <RANKING order="20" place="-1" resultid="4172" />
                    <RANKING order="21" place="-1" resultid="4213" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5819" agemax="9" agemin="9" name="[Maringá] Mirim 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1778" />
                    <RANKING order="2" place="2" resultid="3301" />
                    <RANKING order="3" place="3" resultid="1738" />
                    <RANKING order="4" place="4" resultid="1707" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5820" agemax="10" agemin="10" name="[Maringá] Mirim 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3231" />
                    <RANKING order="2" place="2" resultid="1728" />
                    <RANKING order="3" place="3" resultid="3259" />
                    <RANKING order="4" place="4" resultid="1618" />
                    <RANKING order="5" place="5" resultid="3559" />
                    <RANKING order="6" place="6" resultid="1721" />
                    <RANKING order="7" place="7" resultid="2002" />
                    <RANKING order="8" place="8" resultid="3450" />
                    <RANKING order="9" place="9" resultid="3395" />
                    <RANKING order="10" place="10" resultid="3605" />
                    <RANKING order="11" place="-1" resultid="1733" />
                    <RANKING order="12" place="-1" resultid="3477" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5071" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5072" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5073" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5075" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5076" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5077" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5078" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="5079" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1314" gender="F" number="34" order="6" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5841" agemax="11" agemin="11" name="[Colombo] Petiz 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2466" />
                    <RANKING order="2" place="2" resultid="3959" />
                    <RANKING order="3" place="3" resultid="3279" />
                    <RANKING order="4" place="4" resultid="4242" />
                    <RANKING order="5" place="5" resultid="2968" />
                    <RANKING order="6" place="6" resultid="2438" />
                    <RANKING order="7" place="7" resultid="3380" />
                    <RANKING order="8" place="8" resultid="2550" />
                    <RANKING order="9" place="9" resultid="2487" />
                    <RANKING order="10" place="10" resultid="2445" />
                    <RANKING order="11" place="11" resultid="1855" />
                    <RANKING order="12" place="12" resultid="2051" />
                    <RANKING order="13" place="13" resultid="3938" />
                    <RANKING order="14" place="14" resultid="2501" />
                    <RANKING order="15" place="15" resultid="2620" />
                    <RANKING order="16" place="16" resultid="4007" />
                    <RANKING order="17" place="17" resultid="2646" />
                    <RANKING order="18" place="18" resultid="3979" />
                    <RANKING order="19" place="19" resultid="3700" />
                    <RANKING order="20" place="20" resultid="2716" />
                    <RANKING order="21" place="21" resultid="3366" />
                    <RANKING order="22" place="22" resultid="1908" />
                    <RANKING order="23" place="23" resultid="4184" />
                    <RANKING order="24" place="24" resultid="4055" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5842" agemax="12" agemin="12" name="[Colombo] Petiz 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2515" />
                    <RANKING order="2" place="2" resultid="2389" />
                    <RANKING order="3" place="3" resultid="2473" />
                    <RANKING order="4" place="4" resultid="2335" />
                    <RANKING order="5" place="5" resultid="2382" />
                    <RANKING order="6" place="6" resultid="2328" />
                    <RANKING order="7" place="7" resultid="3952" />
                    <RANKING order="8" place="8" resultid="2947" />
                    <RANKING order="9" place="9" resultid="4111" />
                    <RANKING order="10" place="10" resultid="2709" />
                    <RANKING order="11" place="11" resultid="3925" />
                    <RANKING order="12" place="12" resultid="3462" />
                    <RANKING order="13" place="13" resultid="1848" />
                    <RANKING order="14" place="14" resultid="2410" />
                    <RANKING order="15" place="15" resultid="2459" />
                    <RANKING order="16" place="16" resultid="2375" />
                    <RANKING order="17" place="17" resultid="2081" />
                    <RANKING order="18" place="18" resultid="3784" />
                    <RANKING order="19" place="19" resultid="3353" />
                    <RANKING order="20" place="20" resultid="1882" />
                    <RANKING order="21" place="21" resultid="1375" />
                    <RANKING order="22" place="22" resultid="4144" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5843" agemax="13" agemin="13" name="[Colombo] Infantil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2307" />
                    <RANKING order="2" place="2" resultid="2286" />
                    <RANKING order="3" place="3" resultid="2452" />
                    <RANKING order="4" place="4" resultid="3153" />
                    <RANKING order="5" place="5" resultid="2279" />
                    <RANKING order="6" place="6" resultid="2870" />
                    <RANKING order="7" place="7" resultid="2258" />
                    <RANKING order="8" place="8" resultid="2877" />
                    <RANKING order="9" place="9" resultid="2158" />
                    <RANKING order="10" place="10" resultid="1389" />
                    <RANKING order="11" place="11" resultid="2272" />
                    <RANKING order="12" place="12" resultid="1903" />
                    <RANKING order="13" place="13" resultid="4164" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5844" agemax="14" agemin="14" name="[Colombo] Infantil 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1817" />
                    <RANKING order="2" place="2" resultid="2195" />
                    <RANKING order="3" place="3" resultid="2606" />
                    <RANKING order="4" place="4" resultid="3614" />
                    <RANKING order="5" place="5" resultid="4191" />
                    <RANKING order="6" place="6" resultid="2202" />
                    <RANKING order="7" place="7" resultid="3647" />
                    <RANKING order="8" place="8" resultid="1811" />
                    <RANKING order="9" place="9" resultid="3411" />
                    <RANKING order="10" place="10" resultid="4198" />
                    <RANKING order="11" place="11" resultid="3728" />
                    <RANKING order="12" place="12" resultid="3721" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5845" agemax="15" agemin="15" name="[Colombo] Juvenil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3807" />
                    <RANKING order="2" place="2" resultid="1354" />
                    <RANKING order="3" place="3" resultid="3844" />
                    <RANKING order="4" place="4" resultid="2007" />
                    <RANKING order="5" place="5" resultid="3104" />
                    <RANKING order="6" place="6" resultid="2044" />
                    <RANKING order="7" place="7" resultid="3865" />
                    <RANKING order="8" place="8" resultid="2144" />
                    <RANKING order="9" place="9" resultid="2039" />
                    <RANKING order="10" place="10" resultid="1361" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5846" agemax="-1" agemin="16" name="[Colombo] Juvenil 2/Sênior">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3813" />
                    <RANKING order="2" place="2" resultid="3742" />
                    <RANKING order="3" place="3" resultid="1824" />
                    <RANKING order="4" place="4" resultid="3824" />
                    <RANKING order="5" place="5" resultid="3360" />
                    <RANKING order="6" place="6" resultid="3735" />
                    <RANKING order="7" place="7" resultid="3666" />
                    <RANKING order="8" place="8" resultid="3654" />
                    <RANKING order="9" place="9" resultid="4255" />
                    <RANKING order="10" place="10" resultid="2069" />
                    <RANKING order="11" place="-1" resultid="1843" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5847" agemax="11" agemin="11" name="[Maringá] Petiz 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1680" />
                    <RANKING order="2" place="2" resultid="3314" />
                    <RANKING order="3" place="3" resultid="3265" />
                    <RANKING order="4" place="4" resultid="3244" />
                    <RANKING order="5" place="5" resultid="3251" />
                    <RANKING order="6" place="6" resultid="3132" />
                    <RANKING order="7" place="7" resultid="3216" />
                    <RANKING order="8" place="8" resultid="1610" />
                    <RANKING order="9" place="9" resultid="1570" />
                    <RANKING order="10" place="10" resultid="3490" />
                    <RANKING order="11" place="-1" resultid="1549" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5848" agemax="12" agemin="12" name="[Maringá] Petiz 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3118" />
                    <RANKING order="2" place="2" resultid="3146" />
                    <RANKING order="3" place="3" resultid="1563" />
                    <RANKING order="4" place="4" resultid="3551" />
                    <RANKING order="5" place="5" resultid="1603" />
                    <RANKING order="6" place="6" resultid="3209" />
                    <RANKING order="7" place="7" resultid="3237" />
                    <RANKING order="8" place="8" resultid="3418" />
                    <RANKING order="9" place="9" resultid="3307" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5849" agemax="13" agemin="13" name="[Maringá] Infantil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3286" />
                    <RANKING order="2" place="2" resultid="1500" />
                    <RANKING order="3" place="3" resultid="1975" />
                    <RANKING order="4" place="4" resultid="1493" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5850" agemax="14" agemin="14" name="[Maringá] Infantil 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1936" />
                    <RANKING order="2" place="2" resultid="1963" />
                    <RANKING order="3" place="3" resultid="3571" />
                    <RANKING order="4" place="4" resultid="3181" />
                    <RANKING order="5" place="5" resultid="1486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5851" agemax="15" agemin="15" name="[Maringá] Juvenil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1956" />
                    <RANKING order="2" place="2" resultid="1521" />
                    <RANKING order="3" place="-1" resultid="1528" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5852" agemax="-1" agemin="16" name="[Maringá] Juvenil 2/Sênior">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1949" />
                    <RANKING order="2" place="2" resultid="3525" />
                    <RANKING order="3" place="3" resultid="1514" />
                    <RANKING order="4" place="4" resultid="1767" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5083" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5084" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5085" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5086" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5088" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5089" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5090" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5092" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5093" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="5094" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="5096" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="5097" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="5098" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="5099" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="5100" number="19" order="19" status="OFFICIAL" />
                <HEAT heatid="5101" number="20" order="20" status="OFFICIAL" />
                <HEAT heatid="5102" number="21" order="21" status="OFFICIAL" />
                <HEAT heatid="5103" number="22" order="22" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="4439" gender="F" number="33" order="7" round="FIN" preveventid="1311">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5877" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10173" />
                    <RANKING order="2" place="2" resultid="10174" />
                    <RANKING order="3" place="3" resultid="10175" />
                    <RANKING order="4" place="4" resultid="10179" />
                    <RANKING order="5" place="5" resultid="10177" />
                    <RANKING order="6" place="6" resultid="10178" />
                    <RANKING order="7" place="7" resultid="10039" />
                    <RANKING order="8" place="8" resultid="10040" />
                    <RANKING order="9" place="9" resultid="10043" />
                    <RANKING order="10" place="10" resultid="10042" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5878" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10181" />
                    <RANKING order="2" place="2" resultid="10180" />
                    <RANKING order="3" place="3" resultid="10182" />
                    <RANKING order="4" place="4" resultid="10183" />
                    <RANKING order="5" place="5" resultid="10044" />
                    <RANKING order="6" place="6" resultid="10184" />
                    <RANKING order="7" place="7" resultid="10185" />
                    <RANKING order="8" place="8" resultid="10046" />
                    <RANKING order="9" place="9" resultid="10045" />
                    <RANKING order="10" place="10" resultid="10047" />
                    <RANKING order="11" place="11" resultid="10049" />
                    <RANKING order="12" place="12" resultid="10048" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6048" agegroupid="5877" final="F1" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6049" agegroupid="5877" final="F2" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6050" agegroupid="5878" final="F1" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6051" agegroupid="5878" final="F2" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5804" gender="F" number="34" order="8" round="FIN" preveventid="1314">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5889" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10186" />
                    <RANKING order="2" place="1" resultid="10187" />
                    <RANKING order="3" place="3" resultid="10050" />
                    <RANKING order="4" place="4" resultid="10188" />
                    <RANKING order="5" place="5" resultid="10190" />
                    <RANKING order="6" place="6" resultid="10189" />
                    <RANKING order="7" place="7" resultid="10191" />
                    <RANKING order="8" place="8" resultid="10051" />
                    <RANKING order="9" place="9" resultid="10052" />
                    <RANKING order="10" place="10" resultid="10053" />
                    <RANKING order="11" place="11" resultid="10054" />
                    <RANKING order="12" place="12" resultid="10055" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5890" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10194" />
                    <RANKING order="2" place="2" resultid="10196" />
                    <RANKING order="3" place="3" resultid="10193" />
                    <RANKING order="4" place="4" resultid="10192" />
                    <RANKING order="5" place="5" resultid="10195" />
                    <RANKING order="6" place="6" resultid="10197" />
                    <RANKING order="7" place="7" resultid="10056" />
                    <RANKING order="8" place="8" resultid="10057" />
                    <RANKING order="9" place="9" resultid="10058" />
                    <RANKING order="10" place="10" resultid="10060" />
                    <RANKING order="11" place="11" resultid="10059" />
                    <RANKING order="12" place="12" resultid="10061" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5891" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10200" />
                    <RANKING order="2" place="2" resultid="10201" />
                    <RANKING order="3" place="3" resultid="10199" />
                    <RANKING order="4" place="3" resultid="10202" />
                    <RANKING order="5" place="5" resultid="10198" />
                    <RANKING order="6" place="6" resultid="10203" />
                    <RANKING order="7" place="7" resultid="10066" />
                    <RANKING order="8" place="8" resultid="10064" />
                    <RANKING order="9" place="9" resultid="10062" />
                    <RANKING order="10" place="10" resultid="10065" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5892" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10207" />
                    <RANKING order="2" place="2" resultid="10206" />
                    <RANKING order="3" place="3" resultid="10205" />
                    <RANKING order="4" place="4" resultid="10071" />
                    <RANKING order="5" place="5" resultid="10204" />
                    <RANKING order="6" place="6" resultid="10208" />
                    <RANKING order="7" place="7" resultid="10209" />
                    <RANKING order="8" place="8" resultid="10067" />
                    <RANKING order="9" place="9" resultid="10068" />
                    <RANKING order="10" place="10" resultid="10070" />
                    <RANKING order="11" place="11" resultid="10069" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5893" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10212" />
                    <RANKING order="2" place="2" resultid="10213" />
                    <RANKING order="3" place="3" resultid="10211" />
                    <RANKING order="4" place="4" resultid="10214" />
                    <RANKING order="5" place="5" resultid="10210" />
                    <RANKING order="6" place="6" resultid="10072" />
                    <RANKING order="7" place="7" resultid="10215" />
                    <RANKING order="8" place="8" resultid="10073" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5894" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10218" />
                    <RANKING order="2" place="2" resultid="10219" />
                    <RANKING order="3" place="3" resultid="10217" />
                    <RANKING order="4" place="4" resultid="10220" />
                    <RANKING order="5" place="5" resultid="10076" />
                    <RANKING order="6" place="6" resultid="10216" />
                    <RANKING order="7" place="7" resultid="10222" />
                    <RANKING order="8" place="8" resultid="10075" />
                    <RANKING order="9" place="9" resultid="10074" />
                    <RANKING order="10" place="10" resultid="10077" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6052" agegroupid="5889" final="F1" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6053" agegroupid="5889" final="F2" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6054" agegroupid="5890" final="F1" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6055" agegroupid="5890" final="F2" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6056" agegroupid="5891" final="F1" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6057" agegroupid="5891" final="F2" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6058" agegroupid="5892" final="F1" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6059" agegroupid="5892" final="F2" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6060" agegroupid="5893" final="F1" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6061" agegroupid="5893" final="F2" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6062" agegroupid="5894" final="F1" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="6063" agegroupid="5894" final="F2" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1324" gender="F" number="35" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="8" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1325" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4258" />
                    <RANKING order="2" place="2" resultid="3080" />
                    <RANKING order="3" place="3" resultid="1802" />
                    <RANKING order="4" place="4" resultid="3084" />
                    <RANKING order="5" place="5" resultid="3493" />
                    <RANKING order="6" place="6" resultid="3497" />
                    <RANKING order="7" place="-1" resultid="2120" />
                    <RANKING order="8" place="-1" resultid="2116" />
                    <RANKING order="9" place="-1" resultid="5250" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5122" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5123" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5249" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1326" gender="M" number="36" order="10" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5821" agemax="9" agemin="9" name="[Colombo] Mirim 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2752" />
                    <RANKING order="2" place="2" resultid="2934" />
                    <RANKING order="3" place="3" resultid="2773" />
                    <RANKING order="4" place="4" resultid="4029" />
                    <RANKING order="5" place="5" resultid="3017" />
                    <RANKING order="6" place="6" resultid="2955" />
                    <RANKING order="7" place="7" resultid="1916" />
                    <RANKING order="8" place="8" resultid="2822" />
                    <RANKING order="9" place="9" resultid="3484" />
                    <RANKING order="10" place="10" resultid="4230" />
                    <RANKING order="11" place="11" resultid="2892" />
                    <RANKING order="12" place="12" resultid="2927" />
                    <RANKING order="13" place="13" resultid="3320" />
                    <RANKING order="14" place="14" resultid="2962" />
                    <RANKING order="15" place="-1" resultid="2836" />
                    <RANKING order="16" place="-1" resultid="2899" />
                    <RANKING order="17" place="-1" resultid="2913" />
                    <RANKING order="18" place="-1" resultid="2976" />
                    <RANKING order="19" place="-1" resultid="2989" />
                    <RANKING order="20" place="-1" resultid="2996" />
                    <RANKING order="21" place="-1" resultid="3065" />
                    <RANKING order="22" place="-1" resultid="3071" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5822" agemax="10" agemin="10" name="[Colombo] Mirim 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2600" />
                    <RANKING order="2" place="2" resultid="2696" />
                    <RANKING order="3" place="3" resultid="3974" />
                    <RANKING order="4" place="4" resultid="2586" />
                    <RANKING order="5" place="5" resultid="2689" />
                    <RANKING order="6" place="6" resultid="3024" />
                    <RANKING order="7" place="7" resultid="4077" />
                    <RANKING order="8" place="8" resultid="2885" />
                    <RANKING order="9" place="9" resultid="4098" />
                    <RANKING order="10" place="10" resultid="2661" />
                    <RANKING order="11" place="11" resultid="4105" />
                    <RANKING order="12" place="12" resultid="2593" />
                    <RANKING order="13" place="13" resultid="3994" />
                    <RANKING order="14" place="14" resultid="3967" />
                    <RANKING order="15" place="15" resultid="3429" />
                    <RANKING order="16" place="16" resultid="2668" />
                    <RANKING order="17" place="17" resultid="3078" />
                    <RANKING order="18" place="-1" resultid="1876" />
                    <RANKING order="19" place="-1" resultid="2628" />
                    <RANKING order="20" place="-1" resultid="2635" />
                    <RANKING order="21" place="-1" resultid="2654" />
                    <RANKING order="22" place="-1" resultid="2787" />
                    <RANKING order="23" place="-1" resultid="2808" />
                    <RANKING order="24" place="-1" resultid="4124" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5823" agemax="9" agemin="9" name="[Maringá] Mirim 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1702" />
                    <RANKING order="2" place="2" resultid="1674" />
                    <RANKING order="3" place="3" resultid="3273" />
                    <RANKING order="4" place="4" resultid="3294" />
                    <RANKING order="5" place="5" resultid="1792" />
                    <RANKING order="6" place="-1" resultid="1632" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5824" agemax="10" agemin="10" name="[Maringá] Mirim 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1625" />
                    <RANKING order="2" place="2" resultid="3347" />
                    <RANKING order="3" place="3" resultid="1688" />
                    <RANKING order="4" place="4" resultid="3436" />
                    <RANKING order="5" place="5" resultid="3402" />
                    <RANKING order="6" place="6" resultid="1714" />
                    <RANKING order="7" place="7" resultid="1667" />
                    <RANKING order="8" place="8" resultid="1749" />
                    <RANKING order="9" place="9" resultid="3443" />
                    <RANKING order="10" place="-1" resultid="1785" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5124" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5126" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5127" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5128" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5130" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5131" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5132" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="5133" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="5134" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1329" gender="M" number="37" order="11" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5853" agemax="11" agemin="11" name="[Colombo] Petiz 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3039" />
                    <RANKING order="2" place="2" resultid="1383" />
                    <RANKING order="3" place="3" resultid="4001" />
                    <RANKING order="4" place="4" resultid="2057" />
                    <RANKING order="5" place="5" resultid="2530" />
                    <RANKING order="6" place="6" resultid="4015" />
                    <RANKING order="7" place="7" resultid="2481" />
                    <RANKING order="8" place="7" resultid="2731" />
                    <RANKING order="9" place="9" resultid="4022" />
                    <RANKING order="10" place="10" resultid="2537" />
                    <RANKING order="11" place="11" resultid="2523" />
                    <RANKING order="12" place="12" resultid="2495" />
                    <RANKING order="13" place="13" resultid="3987" />
                    <RANKING order="14" place="14" resultid="3388" />
                    <RANKING order="15" place="15" resultid="4131" />
                    <RANKING order="16" place="16" resultid="3058" />
                    <RANKING order="17" place="17" resultid="3053" />
                    <RANKING order="18" place="18" resultid="3715" />
                    <RANKING order="19" place="-1" resultid="2432" />
                    <RANKING order="20" place="-1" resultid="3326" />
                    <RANKING order="21" place="-1" resultid="2544" />
                    <RANKING order="22" place="-1" resultid="3470" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5854" agemax="12" agemin="12" name="[Colombo] Petiz 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3909" />
                    <RANKING order="2" place="2" resultid="2362" />
                    <RANKING order="3" place="3" resultid="2558" />
                    <RANKING order="4" place="4" resultid="2397" />
                    <RANKING order="5" place="5" resultid="1870" />
                    <RANKING order="6" place="6" resultid="2315" />
                    <RANKING order="7" place="7" resultid="2350" />
                    <RANKING order="8" place="8" resultid="2418" />
                    <RANKING order="9" place="9" resultid="3681" />
                    <RANKING order="10" place="10" resultid="2343" />
                    <RANKING order="11" place="11" resultid="3946" />
                    <RANKING order="12" place="12" resultid="5258" />
                    <RANKING order="13" place="13" resultid="2369" />
                    <RANKING order="14" place="14" resultid="2355" />
                    <RANKING order="15" place="15" resultid="4050" />
                    <RANKING order="16" place="16" resultid="4151" />
                    <RANKING order="17" place="17" resultid="1923" />
                    <RANKING order="18" place="18" resultid="2509" />
                    <RANKING order="19" place="-1" resultid="2404" />
                    <RANKING order="20" place="-1" resultid="2322" />
                    <RANKING order="21" place="-1" resultid="4091" />
                    <RANKING order="22" place="-1" resultid="4236" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5855" agemax="13" agemin="13" name="[Colombo] Infantil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2252" />
                    <RANKING order="2" place="2" resultid="2294" />
                    <RANKING order="3" place="3" resultid="3771" />
                    <RANKING order="4" place="4" resultid="3887" />
                    <RANKING order="5" place="5" resultid="3894" />
                    <RANKING order="6" place="6" resultid="3873" />
                    <RANKING order="7" place="7" resultid="2245" />
                    <RANKING order="8" place="8" resultid="2166" />
                    <RANKING order="9" place="9" resultid="2063" />
                    <RANKING order="10" place="10" resultid="3919" />
                    <RANKING order="11" place="11" resultid="2238" />
                    <RANKING order="12" place="12" resultid="4119" />
                    <RANKING order="13" place="13" resultid="2266" />
                    <RANKING order="14" place="14" resultid="1863" />
                    <RANKING order="15" place="15" resultid="3374" />
                    <RANKING order="16" place="16" resultid="2301" />
                    <RANKING order="17" place="17" resultid="1890" />
                    <RANKING order="18" place="18" resultid="4138" />
                    <RANKING order="19" place="-1" resultid="2173" />
                    <RANKING order="20" place="-1" resultid="2028" />
                    <RANKING order="21" place="-1" resultid="2425" />
                    <RANKING order="22" place="-1" resultid="2565" />
                    <RANKING order="23" place="-1" resultid="3457" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5856" agemax="14" agemin="14" name="[Colombo] Infantil 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3899" />
                    <RANKING order="2" place="2" resultid="2614" />
                    <RANKING order="3" place="3" resultid="2189" />
                    <RANKING order="4" place="4" resultid="2104" />
                    <RANKING order="5" place="5" resultid="10321" />
                    <RANKING order="6" place="6" resultid="4250" />
                    <RANKING order="7" place="7" resultid="2231" />
                    <RANKING order="8" place="8" resultid="4220" />
                    <RANKING order="9" place="9" resultid="2110" />
                    <RANKING order="10" place="10" resultid="2075" />
                    <RANKING order="11" place="11" resultid="3880" />
                    <RANKING order="12" place="12" resultid="2210" />
                    <RANKING order="13" place="13" resultid="3778" />
                    <RANKING order="14" place="14" resultid="2217" />
                    <RANKING order="15" place="15" resultid="4036" />
                    <RANKING order="16" place="16" resultid="4084" />
                    <RANKING order="17" place="-1" resultid="2224" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5857" agemax="15" agemin="15" name="[Colombo] Juvenil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3634" />
                    <RANKING order="2" place="2" resultid="3832" />
                    <RANKING order="3" place="3" resultid="1348" />
                    <RANKING order="4" place="4" resultid="4043" />
                    <RANKING order="5" place="5" resultid="3859" />
                    <RANKING order="6" place="6" resultid="2034" />
                    <RANKING order="7" place="7" resultid="2022" />
                    <RANKING order="8" place="8" resultid="1369" />
                    <RANKING order="9" place="9" resultid="4179" />
                    <RANKING order="10" place="10" resultid="3627" />
                    <RANKING order="11" place="11" resultid="2181" />
                    <RANKING order="12" place="-1" resultid="3839" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5858" agemax="-1" agemin="16" name="[Colombo] Juvenil 2/Sênior">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3641" />
                    <RANKING order="2" place="2" resultid="3333" />
                    <RANKING order="3" place="3" resultid="3792" />
                    <RANKING order="4" place="4" resultid="3708" />
                    <RANKING order="5" place="5" resultid="3687" />
                    <RANKING order="6" place="6" resultid="3799" />
                    <RANKING order="7" place="7" resultid="2138" />
                    <RANKING order="8" place="8" resultid="2152" />
                    <RANKING order="9" place="8" resultid="3694" />
                    <RANKING order="10" place="10" resultid="3852" />
                    <RANKING order="11" place="11" resultid="3620" />
                    <RANKING order="12" place="12" resultid="3820" />
                    <RANKING order="13" place="13" resultid="2015" />
                    <RANKING order="14" place="14" resultid="2089" />
                    <RANKING order="15" place="15" resultid="3340" />
                    <RANKING order="16" place="16" resultid="3660" />
                    <RANKING order="17" place="17" resultid="4206" />
                    <RANKING order="18" place="-1" resultid="3674" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5859" agemax="11" agemin="11" name="[Maringá] Petiz 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1646" />
                    <RANKING order="2" place="2" resultid="1660" />
                    <RANKING order="3" place="3" resultid="1653" />
                    <RANKING order="4" place="4" resultid="1695" />
                    <RANKING order="5" place="5" resultid="1585" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5860" agemax="12" agemin="12" name="[Maringá] Petiz 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1592" />
                    <RANKING order="2" place="2" resultid="1578" />
                    <RANKING order="3" place="3" resultid="3566" />
                    <RANKING order="4" place="4" resultid="1557" />
                    <RANKING order="5" place="5" resultid="3140" />
                    <RANKING order="6" place="6" resultid="3224" />
                    <RANKING order="7" place="7" resultid="1431" />
                    <RANKING order="8" place="8" resultid="3586" />
                    <RANKING order="9" place="9" resultid="1639" />
                    <RANKING order="10" place="10" resultid="1597" />
                    <RANKING order="11" place="11" resultid="3592" />
                    <RANKING order="12" place="-1" resultid="3506" />
                    <RANKING order="13" place="-1" resultid="3598" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5861" agemax="13" agemin="13" name="[Maringá] Infantil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1411" />
                    <RANKING order="2" place="2" resultid="1989" />
                    <RANKING order="3" place="3" resultid="1459" />
                    <RANKING order="4" place="4" resultid="3196" />
                    <RANKING order="5" place="5" resultid="1996" />
                    <RANKING order="6" place="6" resultid="3168" />
                    <RANKING order="7" place="7" resultid="3112" />
                    <RANKING order="8" place="8" resultid="1466" />
                    <RANKING order="9" place="-1" resultid="3175" />
                    <RANKING order="10" place="-1" resultid="3126" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5862" agemax="14" agemin="14" name="[Maringá] Infantil 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3098" />
                    <RANKING order="2" place="2" resultid="1473" />
                    <RANKING order="3" place="3" resultid="3579" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5863" agemax="15" agemin="15" name="[Maringá] Juvenil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1424" />
                    <RANKING order="2" place="2" resultid="3540" />
                    <RANKING order="3" place="3" resultid="1445" />
                    <RANKING order="4" place="4" resultid="3161" />
                    <RANKING order="5" place="5" resultid="3512" />
                    <RANKING order="6" place="-1" resultid="1543" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5864" agemax="-1" agemin="16" name="[Maringá] Juvenil 2/Sênior">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1943" />
                    <RANKING order="2" place="2" resultid="1417" />
                    <RANKING order="3" place="3" resultid="1982" />
                    <RANKING order="4" place="4" resultid="1536" />
                    <RANKING order="5" place="5" resultid="3519" />
                    <RANKING order="6" place="6" resultid="1930" />
                    <RANKING order="7" place="7" resultid="1438" />
                    <RANKING order="8" place="8" resultid="1452" />
                    <RANKING order="9" place="9" resultid="3203" />
                    <RANKING order="10" place="10" resultid="1762" />
                    <RANKING order="11" place="11" resultid="3189" />
                    <RANKING order="12" place="12" resultid="1970" />
                    <RANKING order="13" place="13" resultid="3545" />
                    <RANKING order="14" place="14" resultid="3533" />
                    <RANKING order="15" place="-1" resultid="1755" />
                    <RANKING order="16" place="-1" resultid="1480" />
                    <RANKING order="17" place="-1" resultid="1508" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5137" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5138" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5139" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5140" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5142" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5143" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5144" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5146" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5147" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="5148" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="5150" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="5151" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="5152" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="5154" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="5155" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="5156" number="20" order="20" status="OFFICIAL" />
                <HEAT heatid="5157" number="21" order="21" status="OFFICIAL" />
                <HEAT heatid="5158" number="22" order="22" status="OFFICIAL" />
                <HEAT heatid="5159" number="23" order="23" status="OFFICIAL" />
                <HEAT heatid="5160" number="24" order="24" status="OFFICIAL" />
                <HEAT heatid="5161" number="25" order="25" status="OFFICIAL" />
                <HEAT heatid="5162" number="26" order="26" status="OFFICIAL" />
                <HEAT heatid="5163" number="27" order="27" status="OFFICIAL" />
                <HEAT heatid="5164" number="28" order="28" status="OFFICIAL" />
                <HEAT heatid="5165" number="29" order="29" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="4445" gender="M" number="36" order="12" round="FIN" preveventid="1326">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5879" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10308" />
                    <RANKING order="2" place="2" resultid="10309" />
                    <RANKING order="3" place="3" resultid="10307" />
                    <RANKING order="4" place="4" resultid="10111" />
                    <RANKING order="5" place="5" resultid="10310" />
                    <RANKING order="6" place="6" resultid="10306" />
                    <RANKING order="7" place="7" resultid="10311" />
                    <RANKING order="8" place="8" resultid="10113" />
                    <RANKING order="9" place="9" resultid="10112" />
                    <RANKING order="10" place="10" resultid="10114" />
                    <RANKING order="11" place="11" resultid="10115" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5880" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10116" />
                    <RANKING order="2" place="2" resultid="10314" />
                    <RANKING order="3" place="3" resultid="10315" />
                    <RANKING order="4" place="4" resultid="10312" />
                    <RANKING order="5" place="5" resultid="10313" />
                    <RANKING order="6" place="6" resultid="10316" />
                    <RANKING order="7" place="7" resultid="10317" />
                    <RANKING order="8" place="8" resultid="10117" />
                    <RANKING order="9" place="9" resultid="10119" />
                    <RANKING order="10" place="10" resultid="10118" />
                    <RANKING order="11" place="11" resultid="10120" />
                    <RANKING order="12" place="12" resultid="10121" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6032" agegroupid="5879" final="F1" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6033" agegroupid="5879" final="F2" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6034" agegroupid="5880" final="F1" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6035" agegroupid="5880" final="F2" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5807" gender="M" number="37" order="13" round="FIN" preveventid="1329">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5895" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10269" />
                    <RANKING order="2" place="2" resultid="10270" />
                    <RANKING order="3" place="3" resultid="10271" />
                    <RANKING order="4" place="4" resultid="10122" />
                    <RANKING order="5" place="5" resultid="10267" />
                    <RANKING order="6" place="6" resultid="10272" />
                    <RANKING order="7" place="7" resultid="10123" />
                    <RANKING order="8" place="8" resultid="10125" />
                    <RANKING order="9" place="9" resultid="10124" />
                    <RANKING order="10" place="10" resultid="10126" />
                    <RANKING order="11" place="-1" resultid="10268" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5896" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10276" />
                    <RANKING order="2" place="2" resultid="10275" />
                    <RANKING order="3" place="3" resultid="10274" />
                    <RANKING order="4" place="4" resultid="10277" />
                    <RANKING order="5" place="5" resultid="10127" />
                    <RANKING order="6" place="6" resultid="10273" />
                    <RANKING order="7" place="7" resultid="10128" />
                    <RANKING order="8" place="8" resultid="10129" />
                    <RANKING order="9" place="9" resultid="10278" />
                    <RANKING order="10" place="10" resultid="10130" />
                    <RANKING order="11" place="11" resultid="10131" />
                    <RANKING order="12" place="12" resultid="10132" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5897" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10282" />
                    <RANKING order="2" place="2" resultid="10281" />
                    <RANKING order="3" place="3" resultid="10280" />
                    <RANKING order="4" place="4" resultid="10133" />
                    <RANKING order="5" place="5" resultid="10286" />
                    <RANKING order="6" place="6" resultid="10279" />
                    <RANKING order="7" place="7" resultid="10284" />
                    <RANKING order="8" place="8" resultid="10135" />
                    <RANKING order="9" place="9" resultid="10134" />
                    <RANKING order="10" place="10" resultid="10137" />
                    <RANKING order="11" place="11" resultid="10136" />
                    <RANKING order="12" place="12" resultid="10138" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5898" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10140" />
                    <RANKING order="2" place="2" resultid="10287" />
                    <RANKING order="3" place="3" resultid="10288" />
                    <RANKING order="4" place="4" resultid="10291" />
                    <RANKING order="5" place="5" resultid="10290" />
                    <RANKING order="6" place="6" resultid="10328" />
                    <RANKING order="7" place="7" resultid="10289" />
                    <RANKING order="8" place="8" resultid="10141" />
                    <RANKING order="9" place="-1" resultid="10142" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5899" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10295" />
                    <RANKING order="2" place="2" resultid="10296" />
                    <RANKING order="3" place="3" resultid="10294" />
                    <RANKING order="4" place="4" resultid="10297" />
                    <RANKING order="5" place="5" resultid="10293" />
                    <RANKING order="6" place="6" resultid="10298" />
                    <RANKING order="7" place="7" resultid="10143" />
                    <RANKING order="8" place="8" resultid="10145" />
                    <RANKING order="9" place="9" resultid="10144" />
                    <RANKING order="10" place="10" resultid="10146" />
                    <RANKING order="11" place="11" resultid="10147" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5900" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10149" />
                    <RANKING order="2" place="2" resultid="10148" />
                    <RANKING order="3" place="3" resultid="10151" />
                    <RANKING order="4" place="4" resultid="10150" />
                    <RANKING order="5" place="5" resultid="10152" />
                    <RANKING order="6" place="6" resultid="10301" />
                    <RANKING order="7" place="7" resultid="10153" />
                    <RANKING order="8" place="8" resultid="10300" />
                    <RANKING order="9" place="9" resultid="10303" />
                    <RANKING order="10" place="10" resultid="10299" />
                    <RANKING order="11" place="11" resultid="10305" />
                    <RANKING order="12" place="12" resultid="10304" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6036" agegroupid="5895" final="F1" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="6037" agegroupid="5895" final="F2" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6038" agegroupid="5896" final="F1" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="6039" agegroupid="5896" final="F2" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6040" agegroupid="5897" final="F1" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="6041" agegroupid="5897" final="F2" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6042" agegroupid="5898" final="F1" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="6043" agegroupid="5898" final="F2" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6044" agegroupid="5899" final="F1" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="6045" agegroupid="5899" final="F2" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6046" agegroupid="5900" final="F1" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="6047" agegroupid="5900" final="F2" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1285" gender="M" number="38" order="14" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5825" agemax="9" agemin="9" name="[Colombo] Mirim 1" />
                <AGEGROUP agegroupid="5826" agemax="10" agemin="10" name="[Colombo] Mirim 2" />
                <AGEGROUP agegroupid="5827" agemax="9" agemin="9" name="[Maringá] Mirim 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1701" />
                    <RANKING order="2" place="2" resultid="3272" />
                    <RANKING order="3" place="3" resultid="1673" />
                    <RANKING order="4" place="4" resultid="1791" />
                    <RANKING order="5" place="5" resultid="3293" />
                    <RANKING order="6" place="-1" resultid="1631" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5828" agemax="10" agemin="10" name="[Maringá] Mirim 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1624" />
                    <RANKING order="2" place="2" resultid="1687" />
                    <RANKING order="3" place="3" resultid="1713" />
                    <RANKING order="4" place="4" resultid="3346" />
                    <RANKING order="5" place="5" resultid="3435" />
                    <RANKING order="6" place="6" resultid="3401" />
                    <RANKING order="7" place="7" resultid="1666" />
                    <RANKING order="8" place="8" resultid="1748" />
                    <RANKING order="9" place="9" resultid="3442" />
                    <RANKING order="10" place="-1" resultid="1784" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5192" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="5193" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="5194" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1288" gender="M" number="39" order="15" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5865" agemax="11" agemin="11" name="[Colombo] Petiz 1" />
                <AGEGROUP agegroupid="5866" agemax="12" agemin="12" name="[Colombo] Petiz 2" />
                <AGEGROUP agegroupid="5867" agemax="13" agemin="13" name="[Colombo] Infantil 1" />
                <AGEGROUP agegroupid="5868" agemax="14" agemin="14" name="[Colombo] Infantil 2" />
                <AGEGROUP agegroupid="5869" agemax="15" agemin="15" name="[Colombo] Juvenil 1" />
                <AGEGROUP agegroupid="5870" agemax="-1" agemin="16" name="[Colombo] Juvenil 2/Sênior" />
                <AGEGROUP agegroupid="5871" agemax="11" agemin="11" name="[Maringá] Petiz 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1659" />
                    <RANKING order="2" place="2" resultid="1645" />
                    <RANKING order="3" place="3" resultid="1652" />
                    <RANKING order="4" place="4" resultid="1584" />
                    <RANKING order="5" place="5" resultid="1694" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5872" agemax="12" agemin="12" name="[Maringá] Petiz 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1591" />
                    <RANKING order="2" place="2" resultid="3139" />
                    <RANKING order="3" place="3" resultid="3223" />
                    <RANKING order="4" place="4" resultid="1556" />
                    <RANKING order="5" place="5" resultid="1577" />
                    <RANKING order="6" place="6" resultid="1596" />
                    <RANKING order="7" place="7" resultid="3565" />
                    <RANKING order="8" place="8" resultid="1638" />
                    <RANKING order="9" place="9" resultid="1430" />
                    <RANKING order="10" place="10" resultid="3585" />
                    <RANKING order="11" place="11" resultid="3505" />
                    <RANKING order="12" place="12" resultid="3591" />
                    <RANKING order="13" place="-1" resultid="3597" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5873" agemax="13" agemin="13" name="[Maringá] Infantil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1410" />
                    <RANKING order="2" place="2" resultid="3167" />
                    <RANKING order="3" place="3" resultid="3195" />
                    <RANKING order="4" place="4" resultid="3111" />
                    <RANKING order="5" place="5" resultid="1988" />
                    <RANKING order="6" place="6" resultid="1458" />
                    <RANKING order="7" place="7" resultid="1995" />
                    <RANKING order="8" place="8" resultid="3174" />
                    <RANKING order="9" place="9" resultid="1465" />
                    <RANKING order="10" place="10" resultid="3125" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5874" agemax="14" agemin="14" name="[Maringá] Infantil 2">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3097" />
                    <RANKING order="2" place="2" resultid="1472" />
                    <RANKING order="3" place="3" resultid="3578" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5875" agemax="15" agemin="15" name="[Maringá] Juvenil 1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3539" />
                    <RANKING order="2" place="2" resultid="1423" />
                    <RANKING order="3" place="3" resultid="3511" />
                    <RANKING order="4" place="4" resultid="1444" />
                    <RANKING order="5" place="5" resultid="3160" />
                    <RANKING order="6" place="-1" resultid="1542" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5876" agemax="-1" agemin="16" name="[Maringá] Juvenil 2/Sênior">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1969" />
                    <RANKING order="2" place="2" resultid="1942" />
                    <RANKING order="3" place="3" resultid="1929" />
                    <RANKING order="4" place="4" resultid="3518" />
                    <RANKING order="5" place="5" resultid="1416" />
                    <RANKING order="6" place="6" resultid="1437" />
                    <RANKING order="7" place="7" resultid="1535" />
                    <RANKING order="8" place="8" resultid="1981" />
                    <RANKING order="9" place="9" resultid="3202" />
                    <RANKING order="10" place="10" resultid="1761" />
                    <RANKING order="11" place="11" resultid="3532" />
                    <RANKING order="12" place="12" resultid="1451" />
                    <RANKING order="13" place="13" resultid="3544" />
                    <RANKING order="14" place="14" resultid="3188" />
                    <RANKING order="15" place="15" resultid="1754" />
                    <RANKING order="16" place="-1" resultid="1479" />
                    <RANKING order="17" place="-1" resultid="1507" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5217" number="21" order="21" status="OFFICIAL" />
                <HEAT heatid="5218" number="22" order="22" status="OFFICIAL" />
                <HEAT heatid="5219" number="23" order="23" status="OFFICIAL" />
                <HEAT heatid="5220" number="24" order="24" status="OFFICIAL" />
                <HEAT heatid="5221" number="25" order="25" status="OFFICIAL" />
                <HEAT heatid="5222" number="26" order="26" status="OFFICIAL" />
                <HEAT heatid="5223" number="27" order="27" status="OFFICIAL" />
                <HEAT heatid="5224" number="28" order="28" status="OFFICIAL" />
                <HEAT heatid="5225" number="29" order="29" status="OFFICIAL" />
                <HEAT heatid="5226" number="30" order="30" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="4451" gender="M" number="38" order="16" round="FIN" preveventid="1285">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5881" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10223" />
                    <RANKING order="2" place="2" resultid="10224" />
                    <RANKING order="3" place="3" resultid="10225" />
                    <RANKING order="4" place="4" resultid="10226" />
                    <RANKING order="5" place="5" resultid="10227" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5882" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10229" />
                    <RANKING order="2" place="2" resultid="10230" />
                    <RANKING order="3" place="3" resultid="10232" />
                    <RANKING order="4" place="4" resultid="10233" />
                    <RANKING order="5" place="5" resultid="10231" />
                    <RANKING order="6" place="6" resultid="10234" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6016" agegroupid="5881" final="F1" number="1" order="1" />
                <HEAT heatid="6017" agegroupid="5881" final="F2" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6018" agegroupid="5882" final="F1" number="3" order="3" />
                <HEAT heatid="6019" agegroupid="5882" final="F2" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5810" gender="M" number="39" order="17" round="FIN" preveventid="1288">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5901" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10235" />
                    <RANKING order="2" place="2" resultid="10236" />
                    <RANKING order="3" place="3" resultid="10237" />
                    <RANKING order="4" place="4" resultid="10238" />
                    <RANKING order="5" place="5" resultid="10239" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5902" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10244" />
                    <RANKING order="2" place="2" resultid="10240" />
                    <RANKING order="3" place="3" resultid="10241" />
                    <RANKING order="4" place="4" resultid="10242" />
                    <RANKING order="5" place="5" resultid="10243" />
                    <RANKING order="6" place="6" resultid="10245" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5903" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10246" />
                    <RANKING order="2" place="2" resultid="10247" />
                    <RANKING order="3" place="3" resultid="10248" />
                    <RANKING order="4" place="4" resultid="10250" />
                    <RANKING order="5" place="5" resultid="10249" />
                    <RANKING order="6" place="6" resultid="10251" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5904" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10253" />
                    <RANKING order="2" place="2" resultid="10252" />
                    <RANKING order="3" place="3" resultid="10255" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5905" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10257" />
                    <RANKING order="2" place="2" resultid="10256" />
                    <RANKING order="3" place="3" resultid="10260" />
                    <RANKING order="4" place="4" resultid="10258" />
                    <RANKING order="5" place="5" resultid="10259" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5906" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10261" />
                    <RANKING order="2" place="2" resultid="10262" />
                    <RANKING order="3" place="3" resultid="10263" />
                    <RANKING order="4" place="4" resultid="10264" />
                    <RANKING order="5" place="5" resultid="10266" />
                    <RANKING order="6" place="6" resultid="10265" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6020" agegroupid="5901" final="F1" number="1" order="1" />
                <HEAT heatid="6021" agegroupid="5901" final="F2" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="6022" agegroupid="5902" final="F1" number="3" order="3" />
                <HEAT heatid="6023" agegroupid="5902" final="F2" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="6024" agegroupid="5903" final="F1" number="5" order="5" />
                <HEAT heatid="6025" agegroupid="5903" final="F2" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="6026" agegroupid="5904" final="F1" number="7" order="7" />
                <HEAT heatid="6027" agegroupid="5904" final="F2" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="6028" agegroupid="5905" final="F1" number="9" order="9" />
                <HEAT heatid="6029" agegroupid="5905" final="F2" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="6030" agegroupid="5906" final="F1" number="11" order="11" />
                <HEAT heatid="6031" agegroupid="5906" final="F2" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="10329" gender="M" number="998" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10330" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10445" />
                    <RANKING order="2" place="2" resultid="10382" />
                    <RANKING order="3" place="3" resultid="10461" />
                    <RANKING order="4" place="4" resultid="10522" />
                    <RANKING order="5" place="5" resultid="10444" />
                    <RANKING order="6" place="6" resultid="10471" />
                    <RANKING order="7" place="7" resultid="10539" />
                    <RANKING order="8" place="8" resultid="10482" />
                    <RANKING order="9" place="9" resultid="10451" />
                    <RANKING order="10" place="10" resultid="10455" />
                    <RANKING order="11" place="11" resultid="10448" />
                    <RANKING order="12" place="12" resultid="10454" />
                    <RANKING order="13" place="13" resultid="10456" />
                    <RANKING order="14" place="14" resultid="10457" />
                    <RANKING order="15" place="-1" resultid="10449" />
                    <RANKING order="16" place="-1" resultid="10452" />
                    <RANKING order="17" place="-1" resultid="10453" />
                    <RANKING order="18" place="-1" resultid="10458" />
                    <RANKING order="19" place="-1" resultid="10459" />
                    <RANKING order="20" place="-1" resultid="10460" />
                    <RANKING order="21" place="-1" resultid="10466" />
                    <RANKING order="22" place="-1" resultid="10467" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10331" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10442" />
                    <RANKING order="2" place="2" resultid="10434" />
                    <RANKING order="3" place="3" resultid="10516" />
                    <RANKING order="4" place="4" resultid="10433" />
                    <RANKING order="5" place="5" resultid="10450" />
                    <RANKING order="6" place="6" resultid="10526" />
                    <RANKING order="7" place="7" resultid="10432" />
                    <RANKING order="8" place="8" resultid="10441" />
                    <RANKING order="9" place="9" resultid="10518" />
                    <RANKING order="10" place="10" resultid="10515" />
                    <RANKING order="11" place="11" resultid="10529" />
                    <RANKING order="12" place="12" resultid="10530" />
                    <RANKING order="13" place="13" resultid="10462" />
                    <RANKING order="14" place="14" resultid="10439" />
                    <RANKING order="15" place="15" resultid="10468" />
                    <RANKING order="16" place="-1" resultid="10478" />
                    <RANKING order="17" place="-1" resultid="10380" />
                    <RANKING order="18" place="-1" resultid="10436" />
                    <RANKING order="19" place="-1" resultid="10437" />
                    <RANKING order="20" place="-1" resultid="10438" />
                    <RANKING order="21" place="-1" resultid="10440" />
                    <RANKING order="22" place="-1" resultid="10446" />
                    <RANKING order="23" place="-1" resultid="10447" />
                    <RANKING order="24" place="-1" resultid="10532" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10340" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10341" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10342" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10343" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10344" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10345" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="10332" gender="M" number="999" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10333" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10363" />
                    <RANKING order="2" place="2" resultid="10427" />
                    <RANKING order="3" place="3" resultid="10443" />
                    <RANKING order="4" place="4" resultid="10463" />
                    <RANKING order="5" place="5" resultid="10521" />
                    <RANKING order="6" place="6" resultid="10389" />
                    <RANKING order="7" place="7" resultid="10519" />
                    <RANKING order="8" place="8" resultid="10426" />
                    <RANKING order="9" place="9" resultid="10429" />
                    <RANKING order="10" place="10" resultid="10422" />
                    <RANKING order="11" place="11" resultid="10423" />
                    <RANKING order="12" place="12" resultid="10424" />
                    <RANKING order="13" place="13" resultid="10520" />
                    <RANKING order="14" place="14" resultid="10517" />
                    <RANKING order="15" place="15" resultid="10476" />
                    <RANKING order="16" place="16" resultid="10428" />
                    <RANKING order="17" place="17" resultid="10533" />
                    <RANKING order="18" place="18" resultid="10495" />
                    <RANKING order="19" place="19" resultid="10464" />
                    <RANKING order="20" place="20" resultid="10472" />
                    <RANKING order="21" place="21" resultid="10465" />
                    <RANKING order="22" place="-1" resultid="10481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10334" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10411" />
                    <RANKING order="2" place="2" resultid="10416" />
                    <RANKING order="3" place="3" resultid="10414" />
                    <RANKING order="4" place="4" resultid="10512" />
                    <RANKING order="5" place="5" resultid="10491" />
                    <RANKING order="6" place="6" resultid="10430" />
                    <RANKING order="7" place="7" resultid="10417" />
                    <RANKING order="8" place="8" resultid="10379" />
                    <RANKING order="9" place="9" resultid="10413" />
                    <RANKING order="10" place="10" resultid="10418" />
                    <RANKING order="11" place="11" resultid="10383" />
                    <RANKING order="12" place="12" resultid="10419" />
                    <RANKING order="13" place="13" resultid="10420" />
                    <RANKING order="14" place="14" resultid="10514" />
                    <RANKING order="15" place="15" resultid="10525" />
                    <RANKING order="16" place="16" resultid="10542" />
                    <RANKING order="17" place="17" resultid="10415" />
                    <RANKING order="18" place="18" resultid="10535" />
                    <RANKING order="19" place="19" resultid="10425" />
                    <RANKING order="20" place="-1" resultid="10376" />
                    <RANKING order="21" place="-1" resultid="10377" />
                    <RANKING order="22" place="-1" resultid="10412" />
                    <RANKING order="23" place="-1" resultid="10528" />
                    <RANKING order="24" place="-1" resultid="10540" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10335" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10378" />
                    <RANKING order="2" place="2" resultid="10421" />
                    <RANKING order="3" place="3" resultid="10506" />
                    <RANKING order="4" place="4" resultid="10531" />
                    <RANKING order="5" place="5" resultid="10480" />
                    <RANKING order="6" place="6" resultid="10409" />
                    <RANKING order="7" place="7" resultid="10397" />
                    <RANKING order="8" place="7" resultid="10407" />
                    <RANKING order="9" place="9" resultid="10405" />
                    <RANKING order="10" place="10" resultid="10390" />
                    <RANKING order="11" place="11" resultid="10509" />
                    <RANKING order="12" place="12" resultid="10406" />
                    <RANKING order="13" place="13" resultid="10381" />
                    <RANKING order="14" place="14" resultid="10513" />
                    <RANKING order="15" place="15" resultid="10410" />
                    <RANKING order="16" place="16" resultid="10496" />
                    <RANKING order="17" place="17" resultid="10508" />
                    <RANKING order="18" place="18" resultid="10475" />
                    <RANKING order="19" place="19" resultid="10398" />
                    <RANKING order="20" place="20" resultid="10387" />
                    <RANKING order="21" place="21" resultid="10408" />
                    <RANKING order="22" place="22" resultid="10534" />
                    <RANKING order="23" place="-1" resultid="10431" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10336" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10435" />
                    <RANKING order="2" place="2" resultid="10400" />
                    <RANKING order="3" place="3" resultid="10404" />
                    <RANKING order="4" place="4" resultid="10543" />
                    <RANKING order="5" place="5" resultid="10507" />
                    <RANKING order="6" place="6" resultid="10538" />
                    <RANKING order="7" place="7" resultid="10402" />
                    <RANKING order="8" place="8" resultid="10510" />
                    <RANKING order="9" place="9" resultid="10541" />
                    <RANKING order="10" place="10" resultid="10394" />
                    <RANKING order="11" place="11" resultid="10497" />
                    <RANKING order="12" place="12" resultid="10523" />
                    <RANKING order="13" place="13" resultid="10401" />
                    <RANKING order="14" place="14" resultid="10393" />
                    <RANKING order="15" place="15" resultid="10527" />
                    <RANKING order="16" place="16" resultid="10391" />
                    <RANKING order="17" place="-1" resultid="10403" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10337" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10361" />
                    <RANKING order="2" place="2" resultid="10388" />
                    <RANKING order="3" place="2" resultid="10524" />
                    <RANKING order="4" place="4" resultid="10362" />
                    <RANKING order="5" place="5" resultid="10502" />
                    <RANKING order="6" place="6" resultid="10505" />
                    <RANKING order="7" place="7" resultid="10487" />
                    <RANKING order="8" place="8" resultid="10536" />
                    <RANKING order="9" place="9" resultid="10386" />
                    <RANKING order="10" place="10" resultid="10486" />
                    <RANKING order="11" place="11" resultid="10399" />
                    <RANKING order="12" place="-1" resultid="10503" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10338" agemax="-1" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="10500" />
                    <RANKING order="2" place="2" resultid="10511" />
                    <RANKING order="3" place="3" resultid="10493" />
                    <RANKING order="4" place="4" resultid="10485" />
                    <RANKING order="5" place="5" resultid="10488" />
                    <RANKING order="6" place="6" resultid="10473" />
                    <RANKING order="7" place="7" resultid="10504" />
                    <RANKING order="8" place="8" resultid="10501" />
                    <RANKING order="9" place="9" resultid="10474" />
                    <RANKING order="10" place="10" resultid="10385" />
                    <RANKING order="11" place="11" resultid="10494" />
                    <RANKING order="12" place="12" resultid="10395" />
                    <RANKING order="13" place="13" resultid="10498" />
                    <RANKING order="14" place="14" resultid="10392" />
                    <RANKING order="15" place="15" resultid="10490" />
                    <RANKING order="16" place="16" resultid="10396" />
                    <RANKING order="17" place="17" resultid="10537" />
                    <RANKING order="18" place="18" resultid="10499" />
                    <RANKING order="19" place="19" resultid="10489" />
                    <RANKING order="20" place="20" resultid="10492" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="10346" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="10347" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="10348" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="10349" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="10350" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="10351" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="10352" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="10353" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="10354" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="10355" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="10356" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="10357" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="10358" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="10359" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="10360" number="15" order="15" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1339" gender="M" number="40" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="8" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1340" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4260" />
                    <RANKING order="2" place="2" resultid="10109" />
                    <RANKING order="3" place="3" resultid="3495" />
                    <RANKING order="4" place="4" resultid="3086" />
                    <RANKING order="5" place="5" resultid="3082" />
                    <RANKING order="6" place="-1" resultid="3607" />
                    <RANKING order="7" place="-1" resultid="2122" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5246" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5252" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="1035" nation="BRA" region="PR" clubid="3500" swrid="93778" name="Fundação De Esportes De Campo Mourão" shortname="Fecam">
          <ATHLETES>
            <ATHLETE firstname="Samuel" lastname="Massuda Santos" birthdate="2012-06-09" gender="M" nation="BRA" license="392189" swrid="5603872" athleteid="3560" externalid="392189" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="190" swimtime="00:00:37.80" resultid="3561" heatid="4784" lane="1" />
                <RESULT eventid="1105" points="208" swimtime="00:00:37.27" resultid="3562" heatid="4849" lane="1" entrytime="00:00:40.28" entrycourse="SCM" />
                <RESULT eventid="1249" points="193" swimtime="00:01:23.50" resultid="3563" heatid="4988" lane="5" entrytime="00:01:27.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="221" swimtime="00:01:14.11" resultid="3564" heatid="5015" lane="5" entrytime="00:01:17.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="227" swimtime="00:00:33.01" resultid="3565" heatid="5221" lane="1" entrytime="00:00:33.62" entrycourse="SCM" />
                <RESULT eventid="1329" points="204" swimtime="00:00:42.33" resultid="3566" heatid="5163" lane="1" entrytime="00:00:45.14" entrycourse="SCM" />
                <RESULT eventid="4423" points="191" swimtime="00:00:37.75" resultid="5704" heatid="4795" lane="6" />
                <RESULT eventid="4429" points="206" swimtime="00:00:37.39" resultid="5753" heatid="4855" lane="3" />
                <RESULT eventid="4431" points="223" swimtime="00:00:36.46" resultid="5782" heatid="4865" lane="6" />
                <RESULT eventid="5807" points="223" swimtime="00:00:41.10" resultid="10129" heatid="6039" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaue" lastname="Guilherme Chagas" birthdate="2005-06-29" gender="M" nation="BRA" license="378464" swrid="5603851" athleteid="3541" externalid="378464" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="261" swimtime="00:00:34.01" resultid="3542" heatid="4785" lane="3" />
                <RESULT eventid="1105" points="186" swimtime="00:00:38.68" resultid="3543" heatid="4846" lane="2" />
                <RESULT eventid="1288" points="310" swimtime="00:00:29.78" resultid="3544" heatid="5224" lane="1" entrytime="00:00:28.54" entrycourse="SCM" />
                <RESULT eventid="1329" points="252" swimtime="00:00:39.50" resultid="3545" heatid="5164" lane="2" entrytime="00:00:39.14" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henry" lastname="Sadao Da Silva" birthdate="2012-10-02" gender="M" nation="BRA" license="413907" swrid="5755359" athleteid="3587" externalid="413907" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="69" swimtime="00:00:52.88" resultid="3588" heatid="4783" lane="1" />
                <RESULT eventid="1105" points="69" swimtime="00:00:53.90" resultid="3589" heatid="4846" lane="3" />
                <RESULT eventid="1213" points="71" swimtime="00:02:13.12" resultid="3590" heatid="4957" lane="2" entrytime="00:02:13.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="102" swimtime="00:00:43.10" resultid="3591" heatid="5219" lane="1" entrytime="00:00:43.55" entrycourse="SCM" />
                <RESULT eventid="1329" points="75" swimtime="00:00:59.07" resultid="3592" heatid="5159" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Ferreira Batista" birthdate="2012-03-29" gender="F" nation="BRA" license="385779" swrid="5532525" athleteid="3546" externalid="385779" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="236" swimtime="00:00:39.43" resultid="3547" heatid="4675" lane="3" entrytime="00:00:41.09" entrycourse="SCM" />
                <RESULT eventid="1077" points="220" swimtime="00:00:41.77" resultid="3548" heatid="4727" lane="5" entrytime="00:00:40.97" entrycourse="SCM" />
                <RESULT eventid="1143" points="228" swimtime="00:03:00.52" resultid="3549" heatid="4896" lane="3" entrytime="00:03:00.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                    <SPLIT distance="100" swimtime="00:01:27.64" />
                    <SPLIT distance="150" swimtime="00:02:16.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="238" swimtime="00:01:21.08" resultid="3550" heatid="4938" lane="5" entrytime="00:01:18.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="268" swimtime="00:00:35.55" resultid="3551" heatid="5100" lane="5" entrytime="00:00:35.85" entrycourse="SCM" />
                <RESULT eventid="1301" points="156" swimtime="00:00:52.67" resultid="3552" heatid="5047" lane="1" />
                <RESULT eventid="5804" points="294" swimtime="00:00:34.46" resultid="10059" heatid="6055" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Gomes De Souza" birthdate="2006-01-30" gender="F" nation="BRA" license="308464" swrid="5603844" athleteid="3520" externalid="308464" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="188" swimtime="00:00:42.49" resultid="3521" heatid="4674" lane="2" />
                <RESULT eventid="1077" points="223" swimtime="00:00:41.61" resultid="3522" heatid="4725" lane="6" />
                <RESULT eventid="1129" points="233" swimtime="00:01:41.29" resultid="3523" heatid="4889" lane="4" entrytime="00:01:39.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="212" swimtime="00:03:45.35" resultid="3524" heatid="4923" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.29" />
                    <SPLIT distance="100" swimtime="00:01:42.71" />
                    <SPLIT distance="150" swimtime="00:02:44.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="289" swimtime="00:00:34.67" resultid="3525" heatid="5101" lane="2" entrytime="00:00:33.70" entrycourse="SCM" />
                <RESULT eventid="1301" points="269" swimtime="00:00:43.94" resultid="3526" heatid="5050" lane="3" entrytime="00:00:43.19" entrycourse="SCM" />
                <RESULT eventid="4411" points="183" swimtime="00:00:42.88" resultid="5632" heatid="4689" lane="3" />
                <RESULT eventid="4413" points="178" swimtime="00:00:43.34" resultid="5649" heatid="4695" lane="6" />
                <RESULT eventid="4417" points="240" swimtime="00:00:40.62" resultid="5675" heatid="4740" lane="3" />
                <RESULT eventid="4419" points="245" swimtime="00:00:40.34" resultid="5693" heatid="4746" lane="6" />
                <RESULT eventid="5801" points="264" swimtime="00:00:44.19" resultid="10037" heatid="6077" lane="2" />
                <RESULT eventid="5804" points="291" swimtime="00:00:34.60" resultid="10075" heatid="6063" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Gabrieli Oliveira" birthdate="2010-09-23" gender="F" nation="BRA" license="403428" swrid="5676288" athleteid="3567" externalid="403428" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="229" swimtime="00:00:39.82" resultid="3568" heatid="4675" lane="5" entrytime="00:00:43.78" entrycourse="SCM" />
                <RESULT eventid="1077" points="234" swimtime="00:00:40.96" resultid="3569" heatid="4726" lane="4" entrytime="00:00:43.45" entrycourse="SCM" />
                <RESULT eventid="1189" points="288" swimtime="00:01:16.02" resultid="3570" heatid="4938" lane="2" entrytime="00:01:14.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="309" swimtime="00:00:33.89" resultid="3571" heatid="5101" lane="5" entrytime="00:00:33.97" entrycourse="SCM" />
                <RESULT eventid="1301" points="138" swimtime="00:00:54.82" resultid="3572" heatid="5047" lane="5" />
                <RESULT eventid="4411" points="220" swimtime="00:00:40.36" resultid="5627" heatid="4685" lane="5" />
                <RESULT eventid="4417" points="198" swimtime="00:00:43.32" resultid="5670" heatid="4736" lane="5" />
                <RESULT comment="SW 7.1 - Mais de uma pernada de borboleta antes da primeira pernada de peito após o início ou a virada.  (Horário: 8:58), Após a volta dos 25m." eventid="5801" status="DSQ" swimtime="00:00:53.45" resultid="10031" heatid="6073" lane="5" />
                <RESULT eventid="5804" points="325" swimtime="00:00:33.32" resultid="10069" heatid="6059" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique De Oliveira" birthdate="2009-07-28" gender="M" nation="BRA" license="414505" swrid="5755355" athleteid="3507" externalid="414505" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="376" swimtime="00:00:30.11" resultid="3508" heatid="4790" lane="5" entrytime="00:00:30.36" entrycourse="SCM" />
                <RESULT eventid="1105" points="184" swimtime="00:00:38.82" resultid="3509" heatid="4846" lane="1" />
                <RESULT eventid="1273" points="338" swimtime="00:01:04.32" resultid="3510" heatid="5017" lane="5" entrytime="00:01:04.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="383" swimtime="00:00:27.76" resultid="3511" heatid="5224" lane="5" entrytime="00:00:28.47" entrycourse="SCM" />
                <RESULT eventid="1329" points="238" swimtime="00:00:40.23" resultid="3512" heatid="5157" lane="5" />
                <RESULT eventid="4423" points="346" swimtime="00:00:30.96" resultid="5717" heatid="4801" lane="2" />
                <RESULT eventid="4429" points="191" swimtime="00:00:38.35" resultid="5770" heatid="4861" lane="5" />
                <RESULT eventid="5807" points="220" swimtime="00:00:41.29" resultid="10147" heatid="6045" lane="5" />
                <RESULT eventid="5810" points="369" swimtime="00:00:28.09" resultid="10258" heatid="6029" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Franco Santos" birthdate="2002-01-03" gender="M" nation="BRA" license="290441" swrid="5546064" athleteid="3513" externalid="290441" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="3514" heatid="4791" lane="2" entrytime="00:00:27.37" entrycourse="SCM" />
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="3515" heatid="4843" lane="3" />
                <RESULT eventid="1213" status="DNS" swimtime="00:00:00.00" resultid="3516" heatid="4959" lane="6" entrytime="00:01:17.77" entrycourse="SCM" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="3517" heatid="5018" lane="1" entrytime="00:00:56.96" entrycourse="SCM" />
                <RESULT eventid="1288" points="481" swimtime="00:00:25.72" resultid="3518" heatid="5226" lane="5" entrytime="00:00:25.20" entrycourse="SCM" />
                <RESULT eventid="1329" points="412" swimtime="00:00:33.53" resultid="3519" heatid="5165" lane="5" entrytime="00:00:32.25" entrycourse="SCM" />
                <RESULT eventid="5807" points="418" swimtime="00:00:33.36" resultid="10152" heatid="6047" lane="5" />
                <RESULT eventid="5810" points="500" swimtime="00:00:25.40" resultid="10264" heatid="6031" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Franca Rebollo" birthdate="2012-09-26" gender="M" nation="BRA" license="385780" swrid="5538081" athleteid="3501" externalid="385780" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="100" swimtime="00:00:46.72" resultid="3502" heatid="4786" lane="4" entrytime="00:00:47.55" entrycourse="SCM" />
                <RESULT eventid="1105" points="99" swimtime="00:00:47.68" resultid="3503" heatid="4847" lane="5" entrytime="00:00:50.61" entrycourse="SCM" />
                <RESULT eventid="1273" points="124" swimtime="00:01:29.74" resultid="3504" heatid="5014" lane="4" entrytime="00:01:29.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="120" swimtime="00:00:40.78" resultid="3505" heatid="5219" lane="5" entrytime="00:00:43.18" entrycourse="SCM" />
                <RESULT comment="SW 7.5 - Pés não virados para fora durante a parte propulsora da pernada (fim do ciclo).  (Horário: 10:40)" eventid="1329" status="DSQ" swimtime="00:00:57.65" resultid="3506" heatid="5156" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anthony" lastname="Lira Gordo" birthdate="2012-04-09" gender="M" nation="BRA" license="415261" swrid="5757893" athleteid="3593" externalid="415261" level="MRGA">
              <RESULTS>
                <RESULT comment="SW 8.3 - Movimento alternado das pernas ou pés.  (Horário: 11:44)" eventid="1092" status="DSQ" swimtime="00:00:57.16" resultid="3594" heatid="4782" lane="3" />
                <RESULT eventid="1105" points="72" swimtime="00:00:53.13" resultid="3595" heatid="4844" lane="3" />
                <RESULT eventid="1273" points="108" swimtime="00:01:34.12" resultid="3596" heatid="5013" lane="2" entrytime="00:01:37.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="3597" heatid="5218" lane="5" />
                <RESULT eventid="1329" status="DNS" swimtime="00:00:00.00" resultid="3598" heatid="5161" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stela" lastname="Gouveia" birthdate="2014-02-27" gender="F" nation="BRA" license="415498" swrid="5757891" athleteid="3599" externalid="415498" level="MRGA">
              <RESULTS>
                <RESULT eventid="1061" points="32" swimtime="00:01:16.02" resultid="3600" heatid="4652" lane="3" />
                <RESULT eventid="1074" points="95" swimtime="00:00:55.31" resultid="3601" heatid="4704" lane="4" entrytime="00:00:57.96" entrycourse="SCM" />
                <RESULT eventid="1129" points="67" swimtime="00:02:33.36" resultid="3602" heatid="4888" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="81" swimtime="00:01:56.06" resultid="3603" heatid="4935" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="68" swimtime="00:01:09.33" resultid="3604" heatid="5026" lane="5" />
                <RESULT eventid="1311" points="37" swimtime="00:01:08.79" resultid="3605" heatid="5078" lane="6" entrytime="00:00:51.45" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Stipp Silva" birthdate="2009-12-02" gender="M" nation="BRA" license="378462" swrid="5603918" athleteid="3534" externalid="378462" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="357" swimtime="00:00:30.64" resultid="3535" heatid="4790" lane="6" entrytime="00:00:30.63" entrycourse="SCM" />
                <RESULT eventid="1105" points="268" swimtime="00:00:34.27" resultid="3536" heatid="4846" lane="4" />
                <RESULT eventid="1213" points="360" swimtime="00:01:17.67" resultid="3537" heatid="4958" lane="4" entrytime="00:01:18.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="419" swimtime="00:00:59.92" resultid="3538" heatid="5017" lane="4" entrytime="00:00:59.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="459" swimtime="00:00:26.12" resultid="3539" heatid="5225" lane="4" entrytime="00:00:26.83" entrycourse="SCM" />
                <RESULT eventid="1329" points="361" swimtime="00:00:35.04" resultid="3540" heatid="5164" lane="3" entrytime="00:00:35.86" entrycourse="SCM" />
                <RESULT eventid="4423" points="350" swimtime="00:00:30.86" resultid="5718" heatid="4801" lane="3" />
                <RESULT eventid="4425" points="374" swimtime="00:00:30.17" resultid="5742" heatid="4808" lane="6" />
                <RESULT eventid="4429" points="247" swimtime="00:00:35.21" resultid="5767" heatid="4861" lane="2" />
                <RESULT eventid="4431" points="264" swimtime="00:00:34.44" resultid="5791" heatid="4868" lane="6" />
                <RESULT eventid="5807" points="379" swimtime="00:00:34.47" resultid="10144" heatid="6045" lane="2" />
                <RESULT eventid="5810" points="443" swimtime="00:00:26.43" resultid="10256" heatid="6029" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kenzo" lastname="Kimura" birthdate="2010-04-23" gender="M" nation="BRA" license="403429" swrid="5676289" athleteid="3573" externalid="403429" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="157" swimtime="00:00:40.25" resultid="3574" heatid="4783" lane="5" />
                <RESULT eventid="1105" points="127" swimtime="00:00:43.92" resultid="3575" heatid="4845" lane="4" />
                <RESULT eventid="1227" points="217" swimtime="00:02:45.20" resultid="3576" heatid="5254" lane="2" entrytime="00:02:53.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                    <SPLIT distance="100" swimtime="00:01:15.52" />
                    <SPLIT distance="150" swimtime="00:01:59.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="234" swimtime="00:01:12.71" resultid="3577" heatid="5016" lane="1" entrytime="00:01:12.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="235" swimtime="00:00:32.63" resultid="3578" heatid="5222" lane="6" entrytime="00:00:32.65" entrycourse="SCM" />
                <RESULT eventid="1329" points="208" swimtime="00:00:42.06" resultid="3579" heatid="5163" lane="6" entrytime="00:00:46.96" entrycourse="SCM" />
                <RESULT eventid="4423" points="148" swimtime="00:00:41.10" resultid="5715" heatid="4799" lane="3" />
                <RESULT eventid="4425" points="165" swimtime="00:00:39.58" resultid="5739" heatid="4807" lane="6" />
                <RESULT eventid="4429" points="100" swimtime="00:00:47.50" resultid="5765" heatid="4859" lane="3" />
                <RESULT eventid="4431" points="138" swimtime="00:00:42.77" resultid="5788" heatid="4867" lane="6" />
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 11:10)" eventid="5807" status="DSQ" swimtime="00:00:41.32" resultid="10142" heatid="6043" lane="3" />
                <RESULT eventid="5810" points="238" swimtime="00:00:32.51" resultid="10255" heatid="6027" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Ferreira Batista" birthdate="2014-11-26" gender="F" nation="BRA" license="392160" swrid="5515815" athleteid="3553" externalid="392160" level="MRGA">
              <RESULTS>
                <RESULT eventid="1061" points="78" swimtime="00:00:56.82" resultid="3554" heatid="4653" lane="2" entrytime="00:01:20.79" entrycourse="SCM" />
                <RESULT eventid="1074" points="125" swimtime="00:00:50.38" resultid="3555" heatid="4705" lane="5" entrytime="00:00:52.61" entrycourse="SCM" />
                <RESULT eventid="1165" points="123" swimtime="00:01:50.34" resultid="3556" heatid="4916" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="115" swimtime="00:01:43.08" resultid="3557" heatid="4936" lane="2" entrytime="00:01:50.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="111" swimtime="00:00:58.93" resultid="3558" heatid="5027" lane="2" entrytime="00:01:01.56" entrycourse="SCM" />
                <RESULT eventid="1311" points="156" swimtime="00:00:42.51" resultid="3559" heatid="5078" lane="1" entrytime="00:00:47.35" entrycourse="SCM" />
                <RESULT eventid="4411" points="225" swimtime="00:00:40.03" resultid="5615" heatid="4681" lane="3" />
                <RESULT eventid="4417" points="219" swimtime="00:00:41.83" resultid="5659" heatid="4732" lane="4" />
                <RESULT eventid="4439" points="158" swimtime="00:00:42.40" resultid="10048" heatid="6051" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Eduardo Schork Filho" birthdate="2012-12-28" gender="M" nation="BRA" license="413906" swrid="5755352" athleteid="3580" externalid="413906" level="MRGA">
              <RESULTS>
                <RESULT comment="SW 8.3 - Movimento alternado das pernas ou pés." eventid="1092" status="DSQ" swimtime="00:00:42.58" resultid="3581" heatid="4787" lane="1" entrytime="00:00:45.84" entrycourse="SCM" />
                <RESULT eventid="1105" points="77" swimtime="00:00:51.88" resultid="3582" heatid="4845" lane="1" />
                <RESULT eventid="1213" points="129" swimtime="00:01:49.20" resultid="3583" heatid="4957" lane="4" entrytime="00:01:58.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="130" swimtime="00:01:28.29" resultid="3584" heatid="5014" lane="2" entrytime="00:01:29.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="127" swimtime="00:00:40.03" resultid="3585" heatid="5219" lane="4" entrytime="00:00:42.42" entrycourse="SCM" />
                <RESULT eventid="1329" points="126" swimtime="00:00:49.71" resultid="3586" heatid="5162" lane="4" entrytime="00:00:49.80" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Batinga Ponchielli" birthdate="2007-01-18" gender="M" nation="BRA" license="378461" swrid="5251143" athleteid="3527" externalid="378461" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="186" swimtime="00:00:38.10" resultid="3528" heatid="4785" lane="1" />
                <RESULT eventid="1105" points="244" swimtime="00:00:35.34" resultid="3529" heatid="4849" lane="3" entrytime="00:00:35.13" entrycourse="SCM" />
                <RESULT eventid="1203" points="228" swimtime="00:02:52.79" resultid="3530" heatid="4945" lane="5" entrytime="00:02:53.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                    <SPLIT distance="100" swimtime="00:01:24.76" />
                    <SPLIT distance="150" swimtime="00:02:10.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="231" swimtime="00:01:18.67" resultid="3531" heatid="4988" lane="3" entrytime="00:01:15.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="331" swimtime="00:00:29.12" resultid="3532" heatid="5223" lane="5" entrytime="00:00:29.90" entrycourse="SCM" />
                <RESULT eventid="1329" points="175" swimtime="00:00:44.56" resultid="3533" heatid="5158" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="FECAM/PR &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1115" points="230" swimtime="00:04:52.65" resultid="3606" heatid="5251" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                    <SPLIT distance="100" swimtime="00:01:15.02" />
                    <SPLIT distance="150" swimtime="00:01:53.26" />
                    <SPLIT distance="200" swimtime="00:02:26.35" />
                    <SPLIT distance="250" swimtime="00:02:57.02" />
                    <SPLIT distance="300" swimtime="00:03:36.10" />
                    <SPLIT distance="350" swimtime="00:04:21.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3580" number="1" />
                    <RELAYPOSITION athleteid="3534" number="2" />
                    <RELAYPOSITION athleteid="3560" number="3" />
                    <RELAYPOSITION athleteid="3527" number="4" />
                    <RELAYPOSITION athleteid="3507" number="5" />
                    <RELAYPOSITION athleteid="3541" number="6" />
                    <RELAYPOSITION athleteid="3501" number="7" />
                    <RELAYPOSITION athleteid="3573" number="8" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="SW 10.12 - Os pés perderam contato com a plataforma de partida antes que o colega de equipe anterior tocasse a borda." eventid="1339" status="DSQ" swimtime="00:04:07.29" resultid="3607" heatid="5252" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.16" />
                    <SPLIT distance="100" swimtime="00:01:05.71" />
                    <SPLIT distance="150" swimtime="00:01:33.69" />
                    <SPLIT distance="200" swimtime="00:02:12.63" />
                    <SPLIT distance="250" swimtime="00:02:41.57" />
                    <SPLIT distance="300" swimtime="00:03:09.86" />
                    <SPLIT distance="350" swimtime="00:03:42.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3534" number="1" />
                    <RELAYPOSITION athleteid="3587" number="2" />
                    <RELAYPOSITION athleteid="3527" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="3501" number="4" status="DSQ" />
                    <RELAYPOSITION athleteid="3541" number="5" status="DSQ" />
                    <RELAYPOSITION athleteid="3507" number="6" status="DSQ" />
                    <RELAYPOSITION athleteid="3560" number="7" status="DSQ" />
                    <RELAYPOSITION athleteid="3513" number="8" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="18151" nation="BRA" region="PR" clubid="2174" swrid="95180" name="Clube Uniao Recreativo Palmense" shortname="Clube União">
          <ATHLETES>
            <ATHLETE firstname="Lohan" lastname="Henrique Oliveira" birthdate="2009-03-13" gender="M" nation="BRA" license="410110" swrid="5180392" athleteid="2175" externalid="410110" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="234" swimtime="00:00:35.29" resultid="2176" heatid="4763" lane="1" entrytime="00:00:38.15" entrycourse="SCM" />
                <RESULT eventid="1105" points="188" swimtime="00:00:38.54" resultid="2177" heatid="5253" lane="3" />
                <RESULT eventid="1227" points="265" swimtime="00:02:34.67" resultid="2178" heatid="4966" lane="4" entrytime="00:02:45.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                    <SPLIT distance="100" swimtime="00:01:13.57" />
                    <SPLIT distance="150" swimtime="00:01:55.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="286" swimtime="00:01:08.04" resultid="2179" heatid="5006" lane="1" entrytime="00:01:12.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="239" swimtime="00:00:40.16" resultid="2181" heatid="5154" lane="8" entrytime="00:00:40.35" entrycourse="SCM" />
                <RESULT eventid="10332" points="311" swimtime="00:00:29.75" resultid="10399" heatid="10353" lane="5" entrytime="00:00:32.39" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13068" nation="BRA" region="PR" clubid="3608" swrid="93787" name="Sociedade Morgenau" shortname="Morgenau">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Luiza Melo" birthdate="2015-02-07" gender="F" nation="BRA" license="406717" swrid="5717280" athleteid="3751" externalid="406717" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="95" swimtime="00:00:53.36" resultid="3752" heatid="4649" lane="1" entrytime="00:00:54.98" entrycourse="SCM" />
                <RESULT eventid="1074" points="160" swimtime="00:00:46.44" resultid="3753" heatid="4702" lane="4" entrytime="00:00:44.37" entrycourse="SCM" />
                <RESULT eventid="1165" points="155" swimtime="00:01:42.08" resultid="3754" heatid="4904" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="148" swimtime="00:01:34.90" resultid="3755" heatid="4927" lane="4" entrytime="00:01:34.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="97" swimtime="00:01:01.67" resultid="3756" heatid="5021" lane="8" />
                <RESULT eventid="1311" points="165" swimtime="00:00:41.77" resultid="3757" heatid="5075" lane="1" entrytime="00:00:40.88" entrycourse="SCM" />
                <RESULT eventid="4409" points="97" swimtime="00:00:53.01" resultid="5367" heatid="4655" lane="5" />
                <RESULT eventid="4415" points="157" swimtime="00:00:46.77" resultid="5399" heatid="4706" lane="4" />
                <RESULT eventid="4439" points="161" swimtime="00:00:42.09" resultid="10177" heatid="6048" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Fernanda De Lima" birthdate="2013-09-26" gender="F" nation="BRA" license="378290" swrid="5588693" athleteid="3695" externalid="378290" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="167" swimtime="00:00:44.24" resultid="3696" heatid="4662" lane="3" />
                <RESULT eventid="1077" points="190" swimtime="00:00:43.87" resultid="3697" heatid="4716" lane="6" entrytime="00:00:45.09" entrycourse="SCM" />
                <RESULT eventid="1165" points="188" swimtime="00:01:35.73" resultid="3698" heatid="4911" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="211" swimtime="00:03:05.25" resultid="3699" heatid="4894" lane="2" entrytime="00:03:30.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.32" />
                    <SPLIT distance="100" swimtime="00:01:27.06" />
                    <SPLIT distance="150" swimtime="00:02:18.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="234" swimtime="00:00:37.20" resultid="3700" heatid="5086" lane="3" entrytime="00:00:37.62" entrycourse="SCM" />
                <RESULT eventid="1301" points="139" swimtime="00:00:54.74" resultid="3701" heatid="5040" lane="8" entrytime="00:00:59.75" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolas" lastname="Mingorance Martins" birthdate="2007-10-13" gender="M" nation="BRA" license="393920" swrid="5622295" athleteid="3635" externalid="393920" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="393" swimtime="00:00:29.67" resultid="3636" heatid="4767" lane="3" />
                <RESULT eventid="1105" points="358" swimtime="00:00:31.13" resultid="3637" heatid="4829" lane="4" />
                <RESULT eventid="1227" points="552" swimtime="00:02:01.08" resultid="3638" heatid="4967" lane="3" entrytime="00:02:02.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.30" />
                    <SPLIT distance="100" swimtime="00:00:57.12" />
                    <SPLIT distance="150" swimtime="00:01:28.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="544" swimtime="00:00:54.90" resultid="3639" heatid="5011" lane="5" entrytime="00:00:56.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="384" swimtime="00:00:34.31" resultid="3641" heatid="5154" lane="6" entrytime="00:00:38.22" entrycourse="SCM" />
                <RESULT eventid="4429" points="364" swimtime="00:00:30.94" resultid="5593" heatid="4862" lane="3" />
                <RESULT eventid="4431" points="316" swimtime="00:00:32.44" resultid="5599" heatid="4869" lane="3" />
                <RESULT eventid="5807" points="397" swimtime="00:00:33.92" resultid="10301" heatid="6046" lane="4" />
                <RESULT eventid="10332" points="480" swimtime="00:00:25.74" resultid="10488" heatid="10359" lane="3" entrytime="00:00:25.71" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Kozera Chiarato" birthdate="2010-05-28" gender="M" nation="BRA" license="406722" swrid="5717275" athleteid="3772" externalid="406722" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="321" swimtime="00:00:31.76" resultid="3773" heatid="4778" lane="2" entrytime="00:00:33.97" entrycourse="SCM" />
                <RESULT eventid="1105" points="162" swimtime="00:00:40.53" resultid="3774" heatid="4831" lane="4" />
                <RESULT eventid="1237" points="261" swimtime="00:01:14.75" resultid="3775" heatid="4973" lane="6" entrytime="00:01:18.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="280" swimtime="00:01:08.53" resultid="3776" heatid="5005" lane="4" entrytime="00:01:14.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="202" swimtime="00:00:42.46" resultid="3778" heatid="5152" lane="1" entrytime="00:00:42.48" entrycourse="SCM" />
                <RESULT eventid="10332" points="317" swimtime="00:00:29.56" resultid="10497" heatid="10353" lane="6" entrytime="00:00:32.43" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Tomaz Zmievski" birthdate="2012-09-20" gender="F" nation="BRA" license="406725" swrid="5717300" athleteid="3779" externalid="406725" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="154" swimtime="00:00:45.45" resultid="3780" heatid="4666" lane="4" entrytime="00:00:48.12" entrycourse="SCM" />
                <RESULT eventid="1077" points="196" swimtime="00:00:43.41" resultid="3781" heatid="4714" lane="3" entrytime="00:00:52.62" entrycourse="SCM" />
                <RESULT eventid="1165" points="203" swimtime="00:01:33.25" resultid="3782" heatid="4911" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="248" swimtime="00:02:55.47" resultid="3783" heatid="4894" lane="4" entrytime="00:03:09.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.05" />
                    <SPLIT distance="100" swimtime="00:01:21.28" />
                    <SPLIT distance="150" swimtime="00:02:09.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="266" swimtime="00:00:35.61" resultid="3784" heatid="5086" lane="4" entrytime="00:00:38.00" entrycourse="SCM" />
                <RESULT eventid="1301" points="186" swimtime="00:00:49.66" resultid="3785" heatid="5040" lane="5" entrytime="00:00:56.75" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaylane" lastname="Marques Ferreira" birthdate="2010-03-06" gender="F" nation="BRA" license="391146" swrid="5600211" athleteid="3723" externalid="391146" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="352" swimtime="00:00:34.51" resultid="3724" heatid="4671" lane="1" entrytime="00:00:35.73" entrycourse="SCM" />
                <RESULT eventid="1077" points="203" swimtime="00:00:42.93" resultid="3725" heatid="4712" lane="4" />
                <RESULT eventid="1165" points="175" swimtime="00:01:38.01" resultid="3726" heatid="4907" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="228" swimtime="00:01:28.46" resultid="3727" heatid="4901" lane="5" entrytime="00:01:29.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="292" swimtime="00:00:34.54" resultid="3728" heatid="5090" lane="5" entrytime="00:00:34.66" entrycourse="SCM" />
                <RESULT eventid="1301" points="164" swimtime="00:00:51.77" resultid="3729" heatid="5033" lane="8" />
                <RESULT eventid="4411" points="334" swimtime="00:00:35.13" resultid="5327" heatid="4684" lane="2" />
                <RESULT eventid="4413" points="254" swimtime="00:00:38.47" resultid="5333" heatid="4693" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Nitz Costa" birthdate="2015-02-09" gender="F" nation="BRA" license="397328" swrid="5641773" athleteid="3744" externalid="397328" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="176" swimtime="00:00:43.49" resultid="3745" heatid="4651" lane="5" entrytime="00:00:43.36" entrycourse="SCM" />
                <RESULT eventid="1074" points="196" swimtime="00:00:43.46" resultid="3746" heatid="4702" lane="5" entrytime="00:00:46.36" entrycourse="SCM" />
                <RESULT eventid="1165" points="222" swimtime="00:01:30.54" resultid="3747" heatid="4909" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="246" swimtime="00:01:20.11" resultid="3748" heatid="4928" lane="5" entrytime="00:01:25.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="180" swimtime="00:00:50.17" resultid="3749" heatid="5020" lane="7" />
                <RESULT eventid="1311" points="251" swimtime="00:00:36.34" resultid="3750" heatid="5073" lane="4" entrytime="00:00:43.46" entrycourse="SCM" />
                <RESULT eventid="4409" points="205" swimtime="00:00:41.34" resultid="5364" heatid="4655" lane="2" />
                <RESULT eventid="4415" points="207" swimtime="00:00:42.68" resultid="5396" heatid="4706" lane="1" />
                <RESULT eventid="4433" points="202" swimtime="00:00:48.34" resultid="10081" heatid="5029" lane="3" />
                <RESULT eventid="4439" points="279" swimtime="00:00:35.06" resultid="10173" heatid="6048" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Liz Skowronski" birthdate="2008-01-24" gender="F" nation="BRA" license="358245" swrid="5600202" athleteid="3649" externalid="358245" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="296" swimtime="00:00:36.55" resultid="3650" heatid="4665" lane="6" />
                <RESULT eventid="1077" points="311" swimtime="00:00:37.24" resultid="3651" heatid="4721" lane="4" entrytime="00:00:35.95" entrycourse="SCM" />
                <RESULT eventid="1119" points="341" swimtime="00:02:50.22" resultid="3652" heatid="4876" lane="4" entrytime="00:02:44.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                    <SPLIT distance="100" swimtime="00:01:22.59" />
                    <SPLIT distance="150" swimtime="00:02:06.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="329" swimtime="00:01:19.46" resultid="3653" heatid="4914" lane="1" entrytime="00:01:17.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="355" swimtime="00:00:32.38" resultid="3654" heatid="5083" lane="5" />
                <RESULT eventid="1301" points="258" swimtime="00:00:44.51" resultid="3655" heatid="5033" lane="5" />
                <RESULT eventid="4411" points="277" swimtime="00:00:37.40" resultid="5349" heatid="4688" lane="6" />
                <RESULT eventid="4417" points="321" swimtime="00:00:36.87" resultid="5457" heatid="4739" lane="4" />
                <RESULT eventid="5801" points="256" swimtime="00:00:44.67" resultid="10171" heatid="6076" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Vitor Navarro Zanini" birthdate="2008-06-30" gender="M" nation="BRA" license="369415" swrid="5600273" athleteid="3682" externalid="369415" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="259" swimtime="00:00:34.11" resultid="3683" heatid="4763" lane="5" />
                <RESULT eventid="1105" points="211" swimtime="00:00:37.09" resultid="3684" heatid="4825" lane="2" />
                <RESULT eventid="1213" points="377" swimtime="00:01:16.49" resultid="3685" heatid="4954" lane="6" entrytime="00:01:19.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="361" swimtime="00:00:35.02" resultid="3687" heatid="5155" lane="7" entrytime="00:00:35.40" entrycourse="SCM" />
                <RESULT eventid="5807" points="357" swimtime="00:00:35.15" resultid="10299" heatid="6046" lane="2" />
                <RESULT eventid="10332" points="291" swimtime="00:00:30.42" resultid="10492" heatid="10347" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Rodrigues Galvao" birthdate="2007-04-19" gender="M" nation="BRA" license="376586" swrid="5600247" athleteid="3616" externalid="376586" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="511" swimtime="00:00:27.19" resultid="3617" heatid="4781" lane="4" entrytime="00:00:26.79" entrycourse="SCM" />
                <RESULT eventid="1105" points="380" swimtime="00:00:30.52" resultid="3618" heatid="4823" lane="4" />
                <RESULT eventid="1329" points="293" swimtime="00:00:37.55" resultid="3620" heatid="5144" lane="7" />
                <RESULT eventid="4423" points="505" swimtime="00:00:27.31" resultid="5558" heatid="4802" lane="2" />
                <RESULT eventid="4429" points="370" swimtime="00:00:30.79" resultid="5592" heatid="4862" lane="2" />
                <RESULT eventid="4431" points="309" swimtime="00:00:32.68" resultid="5598" heatid="4869" lane="2" />
                <RESULT eventid="10332" points="481" swimtime="00:00:25.73" resultid="10485" heatid="10360" lane="1" entrytime="00:00:25.45" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduarda" lastname="Azevedo Birsneek" birthdate="2010-03-31" gender="F" nation="BRA" license="391145" swrid="5389427" athleteid="3716" externalid="391145" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="163" swimtime="00:00:44.62" resultid="3717" heatid="4666" lane="2" entrytime="00:00:49.01" entrycourse="SCM" />
                <RESULT eventid="1077" points="186" swimtime="00:00:44.22" resultid="3718" heatid="4716" lane="3" entrytime="00:00:43.18" entrycourse="SCM" />
                <RESULT comment="SW 6.4 - A virada não foi iniciada após a conclusão do movimento de braço, após sair da posição de costas.  (Horário: 16:15), Na volta dos 25m e 75m." eventid="1119" status="DSQ" swimtime="00:03:18.10" resultid="3719" heatid="4876" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.57" />
                    <SPLIT distance="100" swimtime="00:01:37.01" />
                    <SPLIT distance="150" swimtime="00:02:27.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="205" swimtime="00:01:33.09" resultid="3720" heatid="4912" lane="2" entrytime="00:01:36.12" entrycourse="SCM" />
                <RESULT eventid="1314" points="176" swimtime="00:00:40.84" resultid="3721" heatid="5084" lane="4" />
                <RESULT eventid="1301" points="105" swimtime="00:01:00.06" resultid="3722" heatid="5038" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wilson" lastname="Soares Filho" birthdate="2007-12-20" gender="M" nation="BRA" license="414552" swrid="5755379" athleteid="3793" externalid="414552" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="311" swimtime="00:00:32.08" resultid="3794" heatid="4765" lane="3" />
                <RESULT eventid="1105" points="193" swimtime="00:00:38.25" resultid="3795" heatid="4830" lane="4" />
                <RESULT eventid="1227" points="328" swimtime="00:02:24.04" resultid="3796" heatid="4964" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.15" />
                    <SPLIT distance="100" swimtime="00:01:07.17" />
                    <SPLIT distance="150" swimtime="00:01:46.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="324" swimtime="00:01:05.24" resultid="3797" heatid="4998" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="319" swimtime="00:00:36.51" resultid="3799" heatid="5147" lane="1" />
                <RESULT eventid="5807" points="346" swimtime="00:00:35.51" resultid="10305" heatid="6046" lane="7" />
                <RESULT eventid="10332" points="336" swimtime="00:00:28.97" resultid="10499" heatid="10346" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Eduardo Gavinski Alves" birthdate="2012-10-12" gender="M" nation="BRA" license="369324" swrid="5588674" athleteid="3675" externalid="369324" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="228" swimtime="00:00:35.56" resultid="3676" heatid="4775" lane="4" entrytime="00:00:41.09" entrycourse="SCM" />
                <RESULT eventid="1105" points="253" swimtime="00:00:34.95" resultid="3677" heatid="4839" lane="4" entrytime="00:00:34.65" entrycourse="SCM" />
                <RESULT eventid="1203" points="282" swimtime="00:02:40.97" resultid="3678" heatid="4943" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                    <SPLIT distance="100" swimtime="00:01:19.35" />
                    <SPLIT distance="150" swimtime="00:02:01.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="272" swimtime="00:02:33.28" resultid="3679" heatid="4966" lane="2" entrytime="00:02:47.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                    <SPLIT distance="100" swimtime="00:01:12.20" />
                    <SPLIT distance="150" swimtime="00:01:53.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="175" swimtime="00:00:44.55" resultid="3681" heatid="5150" lane="7" entrytime="00:00:51.84" entrycourse="SCM" />
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida." eventid="4429" status="DSQ" swimtime="00:00:34.83" resultid="5521" heatid="4854" lane="2" />
                <RESULT eventid="10332" points="276" swimtime="00:00:30.93" resultid="10491" heatid="10353" lane="4" entrytime="00:00:32.31" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benito" lastname="Alves Sant&apos;Ana" birthdate="2009-06-01" gender="M" nation="BRA" license="376585" swrid="5351951" athleteid="3621" externalid="376585" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="382" swimtime="00:00:29.96" resultid="3622" heatid="4767" lane="6" />
                <RESULT eventid="1105" points="346" swimtime="00:00:31.48" resultid="3623" heatid="4831" lane="5" />
                <RESULT eventid="1203" points="431" swimtime="00:02:19.80" resultid="3624" heatid="4942" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                    <SPLIT distance="100" swimtime="00:01:09.02" />
                    <SPLIT distance="150" swimtime="00:01:45.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1237" points="362" swimtime="00:01:07.01" resultid="3625" heatid="4974" lane="5" entrytime="00:01:10.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="302" swimtime="00:00:37.18" resultid="3627" heatid="5142" lane="4" />
                <RESULT eventid="4429" points="346" swimtime="00:00:31.48" resultid="5589" heatid="4860" lane="5" />
                <RESULT eventid="10332" points="380" swimtime="00:00:27.82" resultid="10486" heatid="10357" lane="5" entrytime="00:00:28.96" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lauren" lastname="Dziura" birthdate="2010-01-11" gender="F" nation="BRA" license="369416" swrid="5588668" athleteid="3642" externalid="369416" level="CLBO">
              <RESULTS>
                <RESULT comment="SW 8.2 - Braços não trazidos para frente simultaneamente sobre (em cima) a água." eventid="1064" status="DSQ" swimtime="00:00:37.88" resultid="3643" heatid="4660" lane="1" />
                <RESULT eventid="1077" points="243" swimtime="00:00:40.42" resultid="3644" heatid="4714" lane="5" />
                <RESULT eventid="1143" points="413" swimtime="00:02:28.10" resultid="3645" heatid="4893" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="380" swimtime="00:01:09.35" resultid="3646" heatid="4926" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="345" swimtime="00:00:32.68" resultid="3647" heatid="5092" lane="6" entrytime="00:00:33.03" entrycourse="SCM" />
                <RESULT eventid="1301" points="260" swimtime="00:00:44.44" resultid="3648" heatid="5034" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Thiago" lastname="Kozera Chiarato" birthdate="2008-01-22" gender="M" nation="BRA" license="406728" swrid="5717276" athleteid="3786" externalid="406728" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="379" swimtime="00:00:30.05" resultid="3787" heatid="4779" lane="2" entrytime="00:00:32.24" entrycourse="SCM" />
                <RESULT eventid="1105" points="265" swimtime="00:00:34.39" resultid="3788" heatid="4832" lane="2" />
                <RESULT eventid="1213" points="378" swimtime="00:01:16.45" resultid="3789" heatid="4948" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="455" swimtime="00:00:58.26" resultid="3790" heatid="5009" lane="2" entrytime="00:01:01.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="372" swimtime="00:00:34.68" resultid="3792" heatid="5154" lane="1" entrytime="00:00:38.80" entrycourse="SCM" />
                <RESULT eventid="5807" points="371" swimtime="00:00:34.72" resultid="10300" heatid="6046" lane="3" />
                <RESULT eventid="10332" points="414" swimtime="00:00:27.04" resultid="10498" heatid="10357" lane="2" entrytime="00:00:28.90" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolas" lastname="Lima" birthdate="2006-12-03" gender="M" nation="BRA" license="366749" swrid="5600201" athleteid="3688" externalid="366749" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="510" swimtime="00:00:27.21" resultid="3689" heatid="4781" lane="2" entrytime="00:00:27.11" entrycourse="SCM" />
                <RESULT eventid="1105" points="257" swimtime="00:00:34.76" resultid="3690" heatid="4823" lane="3" />
                <RESULT eventid="1237" points="500" swimtime="00:01:00.17" resultid="3691" heatid="4974" lane="3" entrytime="00:01:01.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="579" swimtime="00:00:53.77" resultid="3692" heatid="5011" lane="4" entrytime="00:00:54.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="309" swimtime="00:00:36.87" resultid="3694" heatid="5139" lane="4" />
                <RESULT eventid="4423" points="515" swimtime="00:00:27.13" resultid="5559" heatid="4802" lane="3" />
                <RESULT eventid="4425" points="417" swimtime="00:00:29.10" resultid="10318" heatid="4809" lane="3" />
                <RESULT eventid="10332" points="525" swimtime="00:00:24.99" resultid="10493" heatid="10360" lane="4" entrytime="00:00:24.56" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Henrique Opuchkevich" birthdate="2011-02-22" gender="M" nation="BRA" license="406720" swrid="5717273" athleteid="3765" externalid="406720" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="195" swimtime="00:00:37.47" resultid="3766" heatid="4773" lane="5" />
                <RESULT eventid="1105" points="211" swimtime="00:00:37.10" resultid="3767" heatid="4830" lane="3" />
                <RESULT eventid="1227" points="356" swimtime="00:02:20.13" resultid="3768" heatid="4963" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                    <SPLIT distance="100" swimtime="00:01:07.47" />
                    <SPLIT distance="150" swimtime="00:01:44.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="328" swimtime="00:02:54.08" resultid="3769" heatid="4993" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                    <SPLIT distance="100" swimtime="00:01:23.27" />
                    <SPLIT distance="150" swimtime="00:02:09.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="327" swimtime="00:00:36.20" resultid="3771" heatid="5151" lane="4" entrytime="00:00:44.83" entrycourse="SCM" />
                <RESULT eventid="5807" points="330" swimtime="00:00:36.09" resultid="10280" heatid="6040" lane="3" />
                <RESULT eventid="10332" points="280" swimtime="00:00:30.79" resultid="10496" heatid="10351" lane="5" entrytime="00:00:35.36" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Andreis Ramos" birthdate="2007-03-26" gender="M" nation="BRA" license="406719" swrid="5717243" athleteid="3668" externalid="406719" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="375" swimtime="00:00:30.15" resultid="3669" heatid="4778" lane="3" entrytime="00:00:33.28" entrycourse="SCM" />
                <RESULT eventid="1105" points="255" swimtime="00:00:34.85" resultid="3670" heatid="4839" lane="3" entrytime="00:00:34.55" entrycourse="SCM" />
                <RESULT eventid="1237" points="324" swimtime="00:01:09.54" resultid="3671" heatid="4973" lane="3" entrytime="00:01:11.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="375" swimtime="00:01:02.15" resultid="3672" heatid="5008" lane="4" entrytime="00:01:03.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.70" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.5 - Executou uma pernada de borboleta durante o nado." eventid="1329" status="DSQ" swimtime="00:00:36.19" resultid="3674" heatid="5138" lane="2" />
                <RESULT eventid="10332" points="384" swimtime="00:00:27.72" resultid="10490" heatid="10358" lane="6" entrytime="00:00:27.92" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Paes Pereira" birthdate="2013-03-11" gender="M" nation="BRA" license="391137" swrid="5602567" athleteid="3709" externalid="391137" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" status="DSQ" swimtime="00:00:48.10" resultid="3710" heatid="4763" lane="2" />
                <RESULT eventid="1105" points="94" swimtime="00:00:48.52" resultid="3711" heatid="4833" lane="3" />
                <RESULT eventid="1227" points="120" swimtime="00:03:20.91" resultid="3712" heatid="4964" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.32" />
                    <SPLIT distance="100" swimtime="00:01:38.20" />
                    <SPLIT distance="150" swimtime="00:02:32.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="92" swimtime="00:01:46.68" resultid="3713" heatid="4980" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="77" swimtime="00:00:58.56" resultid="3715" heatid="5144" lane="2" />
                <RESULT eventid="10332" points="113" swimtime="00:00:41.60" resultid="10495" heatid="10349" lane="5" entrytime="00:00:42.91" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Luiza Rimbano De Jesus" birthdate="2008-09-02" gender="F" nation="BRA" license="366819" swrid="5653297" athleteid="3737" externalid="366819" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="413" swimtime="00:00:32.73" resultid="3738" heatid="4665" lane="1" />
                <RESULT eventid="1077" points="360" swimtime="00:00:35.49" resultid="3739" heatid="4711" lane="3" />
                <RESULT eventid="1129" points="362" swimtime="00:01:27.46" resultid="3740" heatid="4886" lane="4" entrytime="00:01:26.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="495" swimtime="00:01:03.52" resultid="3741" heatid="4933" lane="4" entrytime="00:01:01.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="488" swimtime="00:00:29.11" resultid="3742" heatid="5097" lane="4" entrytime="00:00:28.40" entrycourse="SCM" />
                <RESULT eventid="1301" points="392" swimtime="00:00:38.76" resultid="3743" heatid="5033" lane="1" />
                <RESULT eventid="4411" points="391" swimtime="00:00:33.32" resultid="5345" heatid="4688" lane="2" />
                <RESULT eventid="4413" points="352" swimtime="00:00:34.50" resultid="5351" heatid="4695" lane="2" />
                <RESULT eventid="4417" points="353" swimtime="00:00:35.72" resultid="5455" heatid="4739" lane="2" />
                <RESULT eventid="4419" points="321" swimtime="00:00:36.84" resultid="5461" heatid="4746" lane="2" />
                <RESULT eventid="5801" points="404" swimtime="00:00:38.35" resultid="10168" heatid="6076" lane="2" />
                <RESULT eventid="5804" points="499" swimtime="00:00:28.89" resultid="10219" heatid="6062" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maryana" lastname="Lemos Carvalho" birthdate="2014-02-10" gender="F" nation="BRA" license="406718" swrid="5717278" athleteid="3758" externalid="406718" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="48" swimtime="00:01:06.68" resultid="3759" heatid="4645" lane="5" />
                <RESULT eventid="1074" points="124" swimtime="00:00:50.59" resultid="3760" heatid="4700" lane="1" entrytime="00:00:52.29" entrycourse="SCM" />
                <RESULT eventid="1165" points="102" swimtime="00:01:57.34" resultid="3761" heatid="4911" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="111" swimtime="00:01:44.48" resultid="3762" heatid="4927" lane="1" entrytime="00:01:41.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="67" swimtime="00:01:09.51" resultid="3763" heatid="5021" lane="7" entrytime="00:01:14.52" entrycourse="SCM" />
                <RESULT eventid="1311" points="162" swimtime="00:00:42.06" resultid="3764" heatid="5072" lane="5" entrytime="00:00:47.59" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kedny" lastname="Correa" birthdate="2004-11-05" gender="M" nation="BRA" license="383858" swrid="5600142" athleteid="3702" externalid="383858" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="419" swimtime="00:00:29.06" resultid="3703" heatid="4780" lane="2" entrytime="00:00:29.60" entrycourse="SCM" />
                <RESULT eventid="1105" points="283" swimtime="00:00:33.67" resultid="3704" heatid="4827" lane="4" />
                <RESULT eventid="1213" points="369" swimtime="00:01:17.04" resultid="3705" heatid="4954" lane="5" entrytime="00:01:16.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="458" swimtime="00:00:58.17" resultid="3706" heatid="4998" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="371" swimtime="00:00:34.70" resultid="3708" heatid="5140" lane="2" />
                <RESULT eventid="4423" points="401" swimtime="00:00:29.48" resultid="5562" heatid="4802" lane="6" />
                <RESULT eventid="5807" points="344" swimtime="00:00:35.58" resultid="10304" heatid="6046" lane="6" />
                <RESULT eventid="10332" points="433" swimtime="00:00:26.64" resultid="10494" heatid="10359" lane="2" entrytime="00:00:26.73" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luana" lastname="Yoshie Kimura" birthdate="2010-07-08" gender="F" nation="BRA" license="391142" swrid="5600277" athleteid="3609" externalid="391142" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="267" swimtime="00:00:37.83" resultid="3610" heatid="4657" lane="3" />
                <RESULT eventid="1077" points="216" swimtime="00:00:42.02" resultid="3611" heatid="4710" lane="5" />
                <RESULT eventid="1129" points="491" swimtime="00:01:19.04" resultid="3612" heatid="4887" lane="3" entrytime="00:01:18.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="440" swimtime="00:02:56.90" resultid="3613" heatid="4922" lane="3" entrytime="00:02:51.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                    <SPLIT distance="100" swimtime="00:01:24.33" />
                    <SPLIT distance="150" swimtime="00:02:11.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="385" swimtime="00:00:31.51" resultid="3614" heatid="5085" lane="8" />
                <RESULT eventid="1301" points="471" swimtime="00:00:36.45" resultid="3615" heatid="5045" lane="3" entrytime="00:00:36.35" entrycourse="SCM" />
                <RESULT eventid="4411" points="295" swimtime="00:00:36.61" resultid="5331" heatid="4684" lane="6" />
                <RESULT eventid="5801" points="488" swimtime="00:00:36.03" resultid="10104" heatid="6072" lane="2" />
                <RESULT eventid="5804" points="389" swimtime="00:00:31.39" resultid="10208" heatid="6058" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Fernanda Pinto" birthdate="2004-09-17" gender="F" nation="BRA" license="391144" swrid="5600157" athleteid="3661" externalid="391144" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="224" swimtime="00:00:40.09" resultid="3662" heatid="4668" lane="1" entrytime="00:00:40.07" entrycourse="SCM" />
                <RESULT eventid="1077" points="248" swimtime="00:00:40.14" resultid="3663" heatid="4717" lane="2" entrytime="00:00:41.66" entrycourse="SCM" />
                <RESULT eventid="1165" points="229" swimtime="00:01:29.68" resultid="3664" heatid="4908" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="333" swimtime="00:01:12.49" resultid="3665" heatid="4930" lane="3" entrytime="00:01:12.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="366" swimtime="00:00:32.04" resultid="3666" heatid="5093" lane="3" entrytime="00:00:31.58" entrycourse="SCM" />
                <RESULT eventid="1301" points="162" swimtime="00:00:51.99" resultid="3667" heatid="5033" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mayara" lastname="Fieber" birthdate="2008-08-20" gender="F" nation="BRA" license="391147" swrid="5600161" athleteid="3730" externalid="391147" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="314" swimtime="00:00:35.86" resultid="3731" heatid="4671" lane="6" entrytime="00:00:35.77" entrycourse="SCM" />
                <RESULT eventid="1077" points="276" swimtime="00:00:38.77" resultid="3732" heatid="4708" lane="2" />
                <RESULT eventid="1153" points="261" swimtime="00:01:24.51" resultid="3733" heatid="4898" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="369" swimtime="00:01:10.00" resultid="3734" heatid="4930" lane="4" entrytime="00:01:13.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="386" swimtime="00:00:31.48" resultid="3735" heatid="5092" lane="3" entrytime="00:00:32.93" entrycourse="SCM" />
                <RESULT eventid="1301" points="342" swimtime="00:00:40.53" resultid="3736" heatid="5042" lane="5" entrytime="00:00:43.76" entrycourse="SCM" />
                <RESULT eventid="4411" points="338" swimtime="00:00:34.97" resultid="5348" heatid="4688" lane="5" />
                <RESULT eventid="4417" points="257" swimtime="00:00:39.68" resultid="5459" heatid="4739" lane="6" />
                <RESULT eventid="5801" points="342" swimtime="00:00:40.55" resultid="10169" heatid="6076" lane="3" />
                <RESULT eventid="5804" points="380" swimtime="00:00:31.64" resultid="10222" heatid="6062" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcus" lastname="Vinicius De Almeida" birthdate="2009-06-16" gender="M" nation="BRA" license="348099" swrid="5600272" athleteid="3628" externalid="348099" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="352" swimtime="00:00:30.79" resultid="3629" heatid="4772" lane="6" />
                <RESULT eventid="1105" points="422" swimtime="00:00:29.46" resultid="3630" heatid="4841" lane="4" entrytime="00:00:30.05" entrycourse="SCM" />
                <RESULT comment="SW 7.1 - Mais de uma pernada de borboleta antes da primeira pernada de peito após o início ou a virada., Na volta dos 25m" eventid="1213" status="DSQ" swimtime="00:01:08.82" resultid="3631" heatid="4954" lane="3" entrytime="00:01:08.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="404" swimtime="00:01:05.33" resultid="3632" heatid="4986" lane="2" entrytime="00:01:05.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="504" swimtime="00:00:31.35" resultid="3634" heatid="5155" lane="4" entrytime="00:00:32.37" entrycourse="SCM" />
                <RESULT eventid="4429" points="427" swimtime="00:00:29.34" resultid="5586" heatid="4860" lane="2" />
                <RESULT eventid="4431" points="387" swimtime="00:00:30.33" resultid="5601" heatid="4868" lane="2" />
                <RESULT eventid="5807" points="520" swimtime="00:00:31.02" resultid="10295" heatid="6044" lane="4" />
                <RESULT eventid="10332" points="413" swimtime="00:00:27.06" resultid="10487" heatid="10346" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Andrianczik Corcini" birthdate="2008-07-19" gender="M" nation="BRA" license="406685" swrid="5736533" athleteid="3656" externalid="406685" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="247" swimtime="00:00:34.65" resultid="3657" heatid="4771" lane="2" />
                <RESULT eventid="1105" points="169" swimtime="00:00:39.93" resultid="3658" heatid="4824" lane="6" />
                <RESULT eventid="1329" points="206" swimtime="00:00:42.21" resultid="3660" heatid="5152" lane="4" entrytime="00:00:40.99" entrycourse="SCM" />
                <RESULT eventid="10332" points="309" swimtime="00:00:29.81" resultid="10489" heatid="10355" lane="3" entrytime="00:00:30.82" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="1007" nation="BRA" region="PR" clubid="3800" swrid="93785" name="Santa Mônica Clube De Campo" shortname="Santa Mônica">
          <ATHLETES>
            <ATHLETE firstname="Bernardo" lastname="Borges Piekarzievicz" birthdate="2013-09-10" gender="M" nation="BRA" license="403142" swrid="5676294" athleteid="4125" externalid="403142" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="67" swimtime="00:00:53.43" resultid="4126" heatid="4763" lane="4" />
                <RESULT eventid="1105" points="103" swimtime="00:00:47.14" resultid="4127" heatid="4834" lane="3" entrytime="00:00:50.55" entrycourse="SCM" />
                <RESULT eventid="1213" status="DNS" swimtime="00:00:00.00" resultid="4128" heatid="4947" lane="6" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="4129" heatid="5001" lane="3" entrytime="00:01:30.16" entrycourse="SCM" />
                <RESULT eventid="1329" points="93" swimtime="00:00:54.97" resultid="4131" heatid="5150" lane="8" entrytime="00:00:52.48" entrycourse="SCM" />
                <RESULT eventid="10332" points="133" swimtime="00:00:39.49" resultid="10533" heatid="10349" lane="4" entrytime="00:00:40.63" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Vicente Lopes" birthdate="2012-03-27" gender="M" nation="BRA" license="415248" swrid="5755344" athleteid="4231" externalid="415248" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="4232" heatid="4769" lane="2" />
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="4233" heatid="4832" lane="6" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="4234" heatid="4997" lane="1" />
                <RESULT eventid="1329" status="DNS" swimtime="00:00:00.00" resultid="4236" heatid="5144" lane="6" />
                <RESULT eventid="10332" status="DNS" swimtime="00:00:00.00" resultid="10540" heatid="10346" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juliana" lastname="Moreira Furtado" birthdate="2011-01-27" gender="F" nation="BRA" license="403783" swrid="5684587" athleteid="4159" externalid="403783" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="141" swimtime="00:00:46.75" resultid="4160" heatid="4661" lane="5" />
                <RESULT eventid="1077" points="200" swimtime="00:00:43.17" resultid="4161" heatid="4708" lane="5" />
                <RESULT eventid="1165" points="209" swimtime="00:01:32.49" resultid="4162" heatid="4912" lane="1" entrytime="00:01:38.32" entrycourse="SCM" />
                <RESULT eventid="1189" points="291" swimtime="00:01:15.80" resultid="4163" heatid="4929" lane="2" entrytime="00:01:19.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="273" swimtime="00:00:35.32" resultid="4164" heatid="5088" lane="6" entrytime="00:00:36.55" entrycourse="SCM" />
                <RESULT eventid="1301" points="132" swimtime="00:00:55.71" resultid="4165" heatid="5032" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Wenceslau Bitencourt" birthdate="2012-02-11" gender="M" nation="BRA" license="377318" swrid="5602591" athleteid="3940" externalid="377318" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="218" swimtime="00:00:36.12" resultid="3941" heatid="4777" lane="1" entrytime="00:00:37.32" entrycourse="SCM" />
                <RESULT eventid="1105" points="183" swimtime="00:00:38.91" resultid="3942" heatid="4836" lane="4" entrytime="00:00:40.07" entrycourse="SCM" />
                <RESULT eventid="1249" points="179" swimtime="00:01:25.73" resultid="3943" heatid="4985" lane="6" entrytime="00:01:27.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="234" swimtime="00:01:12.73" resultid="3944" heatid="4998" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="159" swimtime="00:00:46.03" resultid="3946" heatid="5150" lane="1" entrytime="00:00:52.02" entrycourse="SCM" />
                <RESULT eventid="10332" points="225" swimtime="00:00:33.14" resultid="10514" heatid="10352" lane="3" entrytime="00:00:33.43" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Giuseppe Bulla Lanaro" birthdate="2007-05-22" gender="M" nation="BRA" license="331630" swrid="5600174" athleteid="3808" externalid="331630" level="CLBO">
              <RESULTS>
                <RESULT eventid="1273" points="641" swimtime="00:00:52.00" resultid="3809" heatid="5011" lane="3" entrytime="00:00:52.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10332" points="577" swimtime="00:00:24.21" resultid="10500" heatid="10360" lane="2" entrytime="00:00:24.91" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="Hoffmann Zoschke" birthdate="2015-03-22" gender="M" nation="BRA" license="390917" swrid="5602547" athleteid="4023" externalid="390917" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="132" swimtime="00:00:42.67" resultid="4024" heatid="4755" lane="2" entrytime="00:00:46.92" entrycourse="SCM" />
                <RESULT eventid="1102" points="110" swimtime="00:00:46.04" resultid="4025" heatid="4810" lane="5" />
                <RESULT eventid="1213" points="113" swimtime="00:01:54.32" resultid="4026" heatid="4949" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="176" swimtime="00:01:19.92" resultid="4027" heatid="5004" lane="3" entrytime="00:01:19.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="114" swimtime="00:00:51.40" resultid="4029" heatid="5128" lane="7" entrytime="00:00:56.60" entrycourse="SCM" />
                <RESULT eventid="4421" points="148" swimtime="00:00:41.04" resultid="5464" heatid="4760" lane="2" />
                <RESULT eventid="4427" points="110" swimtime="00:00:46.03" resultid="5502" heatid="4821" lane="4" />
                <RESULT eventid="4445" points="122" swimtime="00:00:50.23" resultid="10310" heatid="6032" lane="6" />
                <RESULT eventid="10329" points="158" swimtime="00:00:37.25" resultid="10522" heatid="10344" lane="3" entrytime="00:00:36.35" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="De Siqueira Machado" birthdate="2012-05-25" gender="F" nation="BRA" license="377312" swrid="5588649" athleteid="3920" externalid="377312" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="291" swimtime="00:00:36.76" resultid="3921" heatid="4669" lane="4" entrytime="00:00:38.21" entrycourse="SCM" />
                <RESULT eventid="1077" points="255" swimtime="00:00:39.81" resultid="3922" heatid="4720" lane="2" entrytime="00:00:37.77" entrycourse="SCM" />
                <RESULT eventid="1119" points="213" swimtime="00:03:19.05" resultid="3923" heatid="4875" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.09" />
                    <SPLIT distance="100" swimtime="00:01:35.70" />
                    <SPLIT distance="150" swimtime="00:02:27.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="310" swimtime="00:01:14.19" resultid="3924" heatid="4930" lane="1" entrytime="00:01:14.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="359" swimtime="00:00:32.25" resultid="3925" heatid="5094" lane="7" entrytime="00:00:30.76" entrycourse="SCM" />
                <RESULT eventid="1301" points="292" swimtime="00:00:42.75" resultid="3926" heatid="5042" lane="3" entrytime="00:00:42.93" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Marini" birthdate="2014-04-09" gender="M" nation="BRA" license="382247" swrid="5684582" athleteid="3961" externalid="382247" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="106" swimtime="00:00:45.84" resultid="3962" heatid="4755" lane="1" entrytime="00:00:48.08" entrycourse="SCM" />
                <RESULT eventid="1102" points="119" swimtime="00:00:44.84" resultid="3963" heatid="4815" lane="1" entrytime="00:00:50.75" entrycourse="SCM" />
                <RESULT eventid="1249" points="120" swimtime="00:01:37.84" resultid="3964" heatid="4979" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="122" swimtime="00:01:30.29" resultid="3965" heatid="5003" lane="2" entrytime="00:01:26.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="91" swimtime="00:00:55.36" resultid="3967" heatid="5128" lane="4" entrytime="00:01:01.79" entrycourse="SCM" />
                <RESULT eventid="10329" points="136" swimtime="00:00:39.13" resultid="10515" heatid="10343" lane="3" entrytime="00:00:39.78" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Zanardi" birthdate="2008-10-02" gender="F" nation="BRA" license="398572" swrid="5757089" athleteid="4251" externalid="398572" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="239" swimtime="00:00:39.24" resultid="4252" heatid="4661" lane="1" />
                <RESULT eventid="1077" points="220" swimtime="00:00:41.77" resultid="4253" heatid="4712" lane="1" />
                <RESULT eventid="1165" points="207" swimtime="00:01:32.66" resultid="4254" heatid="4910" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="284" swimtime="00:00:34.87" resultid="4255" heatid="5090" lane="1" entrytime="00:00:34.86" entrycourse="SCM" />
                <RESULT eventid="1301" points="227" swimtime="00:00:46.46" resultid="4256" heatid="5041" lane="4" entrytime="00:00:46.61" entrycourse="SCM" />
                <RESULT eventid="5801" points="197" swimtime="00:00:48.74" resultid="10172" heatid="6076" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Cardim Martins" birthdate="2010-09-01" gender="F" nation="BRA" license="390920" swrid="5600130" athleteid="4193" externalid="390920" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="237" swimtime="00:00:39.36" resultid="4194" heatid="4668" lane="6" entrytime="00:00:40.47" entrycourse="SCM" />
                <RESULT eventid="1077" points="280" swimtime="00:00:38.56" resultid="4195" heatid="4718" lane="5" entrytime="00:00:40.70" entrycourse="SCM" />
                <RESULT eventid="1119" points="328" swimtime="00:02:52.30" resultid="4196" heatid="4875" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.91" />
                    <SPLIT distance="100" swimtime="00:01:24.28" />
                    <SPLIT distance="150" swimtime="00:02:09.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="309" swimtime="00:01:21.19" resultid="4197" heatid="4910" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="296" swimtime="00:00:34.40" resultid="4198" heatid="5089" lane="8" entrytime="00:00:36.35" entrycourse="SCM" />
                <RESULT eventid="1301" points="216" swimtime="00:00:47.28" resultid="4199" heatid="5033" lane="4" />
                <RESULT eventid="4417" points="284" swimtime="00:00:38.41" resultid="5439" heatid="4735" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helenna" lastname="Banzatto Silva" birthdate="2013-07-11" gender="F" nation="BRA" license="393210" swrid="5616439" athleteid="4051" externalid="393210" level="CLBO">
              <RESULTS>
                <RESULT comment="SW 8.3 - Movimento alternado das pernas ou pés." eventid="1064" status="DSQ" swimtime="00:01:10.21" resultid="4052" heatid="4661" lane="2" />
                <RESULT eventid="1077" points="67" swimtime="00:01:01.93" resultid="4053" heatid="4714" lane="2" entrytime="00:01:13.25" entrycourse="SCM" />
                <RESULT eventid="1129" points="154" swimtime="00:01:56.10" resultid="4054" heatid="4884" lane="3" entrytime="00:01:58.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="89" swimtime="00:00:51.28" resultid="4055" heatid="5085" lane="4" entrytime="00:00:52.64" entrycourse="SCM" />
                <RESULT comment="SW 7.1 - Mais de uma pernada de borboleta antes da primeira pernada de peito após o início ou a virada., Após a volta dsos 25m." eventid="1301" status="DSQ" swimtime="00:00:54.47" resultid="4056" heatid="5040" lane="1" entrytime="00:00:55.29" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otavio" lastname="Andrade Guarido" birthdate="2014-05-17" gender="M" nation="BRA" license="400031" swrid="5652873" athleteid="4092" externalid="400031" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="72" swimtime="00:00:52.25" resultid="4093" heatid="4749" lane="4" />
                <RESULT eventid="1102" points="92" swimtime="00:00:48.89" resultid="4094" heatid="4814" lane="2" entrytime="00:00:54.39" entrycourse="SCM" />
                <RESULT eventid="1213" points="116" swimtime="00:01:53.23" resultid="4095" heatid="4949" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="113" swimtime="00:01:32.69" resultid="4096" heatid="5000" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="103" swimtime="00:00:53.11" resultid="4098" heatid="5131" lane="8" entrytime="00:00:53.22" entrycourse="SCM" />
                <RESULT eventid="10329" points="135" swimtime="00:00:39.21" resultid="10529" heatid="10344" lane="1" entrytime="00:00:39.16" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Inoue Kuroda" birthdate="2009-04-18" gender="M" nation="BRA" license="324700" swrid="5600190" athleteid="3833" externalid="324700" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="3834" heatid="4768" lane="3" />
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="3835" heatid="4841" lane="5" entrytime="00:00:30.85" entrycourse="SCM" />
                <RESULT eventid="1227" status="DNS" swimtime="00:00:00.00" resultid="3836" heatid="4967" lane="4" entrytime="00:02:04.17" entrycourse="SCM" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="3837" heatid="5010" lane="3" entrytime="00:00:58.06" entrycourse="SCM" />
                <RESULT eventid="1329" status="DNS" swimtime="00:00:00.00" resultid="3839" heatid="5140" lane="8" />
                <RESULT eventid="10332" status="DNS" swimtime="00:00:00.00" resultid="10503" heatid="10359" lane="6" entrytime="00:00:26.61" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Gouvea" birthdate="2013-04-19" gender="M" nation="BRA" license="387378" swrid="5588729" athleteid="3995" externalid="387378" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="129" swimtime="00:00:42.98" resultid="3996" heatid="4774" lane="3" entrytime="00:00:49.28" entrycourse="SCM" />
                <RESULT eventid="1105" points="172" swimtime="00:00:39.69" resultid="3997" heatid="4829" lane="2" />
                <RESULT eventid="1213" points="190" swimtime="00:01:36.03" resultid="3998" heatid="4952" lane="5" entrytime="00:01:36.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="188" swimtime="00:03:29.60" resultid="3999" heatid="4992" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.14" />
                    <SPLIT distance="100" swimtime="00:01:40.85" />
                    <SPLIT distance="150" swimtime="00:02:35.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="209" swimtime="00:00:42.01" resultid="4001" heatid="5151" lane="1" entrytime="00:00:45.35" entrycourse="SCM" />
                <RESULT eventid="4429" points="182" swimtime="00:00:38.98" resultid="5514" heatid="4852" lane="4" />
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida." eventid="5807" status="DSQ" swimtime="00:00:42.91" resultid="10268" heatid="6036" lane="3" />
                <RESULT eventid="10332" points="230" swimtime="00:00:32.90" resultid="10519" heatid="10352" lane="5" entrytime="00:00:34.63" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Strapasson" birthdate="2012-03-01" gender="M" nation="BRA" license="371377" swrid="5602585" athleteid="3903" externalid="371377" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="239" swimtime="00:00:35.00" resultid="3904" heatid="4768" lane="5" />
                <RESULT eventid="1105" points="165" swimtime="00:00:40.31" resultid="3905" heatid="4823" lane="2" />
                <RESULT eventid="1263" points="281" swimtime="00:03:03.33" resultid="3906" heatid="4992" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.64" />
                    <SPLIT distance="100" swimtime="00:01:26.30" />
                    <SPLIT distance="150" swimtime="00:02:15.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="310" swimtime="00:01:06.19" resultid="3907" heatid="5007" lane="3" entrytime="00:01:06.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="299" swimtime="00:00:37.29" resultid="3909" heatid="5154" lane="7" entrytime="00:00:39.17" entrycourse="SCM" />
                <RESULT eventid="4425" points="226" swimtime="00:00:35.67" resultid="5605" heatid="4805" lane="3" />
                <RESULT eventid="5807" points="291" swimtime="00:00:37.61" resultid="10275" heatid="6038" lane="4" />
                <RESULT eventid="4423" points="255" swimtime="00:00:34.28" resultid="10324" heatid="4794" lane="5" />
                <RESULT eventid="10332" points="310" swimtime="00:00:29.76" resultid="10512" heatid="10356" lane="5" entrytime="00:00:29.78" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Vianna" birthdate="2011-01-31" gender="M" nation="BRA" license="371380" swrid="5588947" athleteid="3910" externalid="371380" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="301" swimtime="00:00:32.44" resultid="3911" heatid="4764" lane="3" />
                <RESULT eventid="1105" points="221" swimtime="00:00:36.53" resultid="3912" heatid="4826" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Bello Costa Lange" birthdate="2010-09-13" gender="M" nation="BRA" license="367152" swrid="5588547" athleteid="3895" externalid="367152" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="378" swimtime="00:00:30.06" resultid="3896" heatid="4779" lane="1" entrytime="00:00:32.36" entrycourse="SCM" />
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="3897" heatid="4824" lane="5" />
                <RESULT eventid="1329" points="360" swimtime="00:00:35.05" resultid="3899" heatid="5144" lane="4" />
                <RESULT eventid="4423" points="396" swimtime="00:00:29.61" resultid="5541" heatid="4798" lane="4" />
                <RESULT eventid="5807" points="362" swimtime="00:00:34.99" resultid="10288" heatid="6042" lane="4" />
                <RESULT eventid="4425" points="361" swimtime="00:00:30.53" resultid="10325" heatid="4807" lane="2" />
                <RESULT eventid="10332" points="356" swimtime="00:00:28.43" resultid="10510" heatid="10357" lane="7" entrytime="00:00:29.79" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Marques Machado" birthdate="2010-02-17" gender="M" nation="BRA" license="390918" swrid="5600212" athleteid="4030" externalid="390918" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="324" swimtime="00:00:31.66" resultid="4031" heatid="4764" lane="6" />
                <RESULT eventid="1105" points="188" swimtime="00:00:38.53" resultid="4032" heatid="4825" lane="6" />
                <RESULT eventid="1227" points="377" swimtime="00:02:17.47" resultid="4033" heatid="4964" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                    <SPLIT distance="100" swimtime="00:01:06.74" />
                    <SPLIT distance="150" swimtime="00:01:42.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1237" points="273" swimtime="00:01:13.63" resultid="4034" heatid="4969" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="193" swimtime="00:00:43.13" resultid="4036" heatid="5138" lane="7" />
                <RESULT eventid="4423" points="311" swimtime="00:00:32.07" resultid="5543" heatid="4798" lane="6" />
                <RESULT eventid="10332" points="314" swimtime="00:00:29.65" resultid="10523" heatid="10348" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Camily Moraes" birthdate="2014-07-13" gender="F" nation="BRA" license="397159" swrid="5641755" athleteid="4064" externalid="397159" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="107" swimtime="00:00:51.28" resultid="4065" heatid="4645" lane="1" />
                <RESULT eventid="1074" points="170" swimtime="00:00:45.55" resultid="4066" heatid="4701" lane="3" entrytime="00:00:48.12" entrycourse="SCM" />
                <RESULT eventid="1129" points="195" swimtime="00:01:47.49" resultid="4067" heatid="4879" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="158" swimtime="00:01:41.42" resultid="4068" heatid="4907" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="166" swimtime="00:00:51.61" resultid="4069" heatid="5023" lane="3" entrytime="00:01:03.23" entrycourse="SCM" />
                <RESULT eventid="1311" points="200" swimtime="00:00:39.17" resultid="4070" heatid="5076" lane="6" entrytime="00:00:39.56" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Leticia Durat" birthdate="2008-02-09" gender="F" nation="BRA" license="331636" swrid="5600200" athleteid="3821" externalid="331636" level="CLBO">
              <RESULTS>
                <RESULT eventid="1129" points="343" swimtime="00:01:29.07" resultid="3822" heatid="4881" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="316" swimtime="00:03:17.43" resultid="3823" heatid="4921" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.94" />
                    <SPLIT distance="100" swimtime="00:01:34.13" />
                    <SPLIT distance="150" swimtime="00:02:24.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="399" swimtime="00:00:31.14" resultid="3824" heatid="5094" lane="4" entrytime="00:00:30.89" entrycourse="SCM" />
                <RESULT eventid="1301" points="335" swimtime="00:00:40.82" resultid="3825" heatid="5036" lane="2" />
                <RESULT eventid="5801" points="351" swimtime="00:00:40.21" resultid="10170" heatid="6076" lane="4" />
                <RESULT eventid="5804" points="392" swimtime="00:00:31.32" resultid="10220" heatid="6062" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Blansky Hagebock" birthdate="2008-08-15" gender="M" nation="BRA" license="339123" swrid="5455418" athleteid="3846" externalid="339123" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="444" swimtime="00:00:28.49" resultid="3847" heatid="4780" lane="4" entrytime="00:00:29.00" entrycourse="SCM" />
                <RESULT eventid="1105" points="299" swimtime="00:00:33.05" resultid="3848" heatid="4834" lane="6" />
                <RESULT eventid="1227" points="498" swimtime="00:02:05.31" resultid="3849" heatid="4967" lane="5" entrytime="00:02:09.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.84" />
                    <SPLIT distance="100" swimtime="00:01:00.21" />
                    <SPLIT distance="150" swimtime="00:01:33.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="561" swimtime="00:00:54.35" resultid="3850" heatid="5011" lane="2" entrytime="00:00:55.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="293" swimtime="00:00:37.53" resultid="3852" heatid="5137" lane="6" />
                <RESULT eventid="4423" points="388" swimtime="00:00:29.82" resultid="5561" heatid="4802" lane="5" />
                <RESULT eventid="4429" points="282" swimtime="00:00:33.68" resultid="5596" heatid="4862" lane="6" />
                <RESULT eventid="10332" points="469" swimtime="00:00:25.93" resultid="10504" heatid="10359" lane="4" entrytime="00:00:26.07" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Faustino Canjerana" birthdate="2013-09-27" gender="F" nation="BRA" license="416735" swrid="5756905" athleteid="4237" externalid="416735" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="306" swimtime="00:00:36.17" resultid="4238" heatid="4658" lane="2" />
                <RESULT eventid="1077" points="193" swimtime="00:00:43.69" resultid="4239" heatid="4713" lane="1" />
                <RESULT eventid="1143" points="312" swimtime="00:02:42.60" resultid="4240" heatid="4894" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.68" />
                    <SPLIT distance="100" swimtime="00:01:19.59" />
                    <SPLIT distance="150" swimtime="00:02:03.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="342" swimtime="00:01:11.83" resultid="4241" heatid="4926" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="354" swimtime="00:00:32.39" resultid="4242" heatid="5084" lane="8" />
                <RESULT eventid="1301" points="225" swimtime="00:00:46.60" resultid="4243" heatid="5034" lane="7" />
                <RESULT eventid="4413" points="258" swimtime="00:00:38.26" resultid="5377" heatid="4690" lane="3" />
                <RESULT eventid="4411" points="322" swimtime="00:00:35.56" resultid="5383" heatid="4678" lane="3" />
                <RESULT eventid="5804" points="345" swimtime="00:00:32.67" resultid="10189" heatid="6052" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Larissa" lastname="Araujo Felix" birthdate="2010-05-27" gender="F" nation="BRA" license="393157" swrid="5622260" athleteid="4186" externalid="393157" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="286" swimtime="00:00:36.97" resultid="4187" heatid="4665" lane="2" />
                <RESULT eventid="1077" points="326" swimtime="00:00:36.68" resultid="4188" heatid="4713" lane="2" />
                <RESULT eventid="1165" points="293" swimtime="00:01:22.57" resultid="4189" heatid="4908" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="355" swimtime="00:01:10.92" resultid="4190" heatid="4926" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="362" swimtime="00:00:32.16" resultid="4191" heatid="5089" lane="4" entrytime="00:00:35.16" entrycourse="SCM" />
                <RESULT eventid="1301" points="177" swimtime="00:00:50.49" resultid="4192" heatid="5037" lane="8" />
                <RESULT eventid="4411" points="314" swimtime="00:00:35.84" resultid="5330" heatid="4684" lane="5" />
                <RESULT eventid="4417" points="318" swimtime="00:00:36.99" resultid="5437" heatid="4735" lane="2" />
                <RESULT eventid="4419" points="265" swimtime="00:00:39.31" resultid="5443" heatid="4744" lane="2" />
                <RESULT eventid="5804" points="403" swimtime="00:00:31.04" resultid="10204" heatid="6058" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexandre" lastname="Celli Schneider" birthdate="2011-02-21" gender="M" nation="BRA" license="367055" swrid="5588587" athleteid="3867" externalid="367055" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="358" swimtime="00:00:30.63" resultid="3868" heatid="4764" lane="5" />
                <RESULT eventid="1105" points="302" swimtime="00:00:32.94" resultid="3869" heatid="4840" lane="5" entrytime="00:00:33.78" entrycourse="SCM" />
                <RESULT eventid="1203" points="343" swimtime="00:02:30.81" resultid="3870" heatid="4943" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                    <SPLIT distance="100" swimtime="00:01:13.53" />
                    <SPLIT distance="150" swimtime="00:01:53.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1237" points="326" swimtime="00:01:09.36" resultid="3871" heatid="4973" lane="2" entrytime="00:01:14.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="279" swimtime="00:00:38.18" resultid="3873" heatid="5139" lane="5" />
                <RESULT eventid="4423" points="366" swimtime="00:00:30.38" resultid="5531" heatid="4796" lane="3" />
                <RESULT eventid="4425" points="324" swimtime="00:00:31.64" resultid="5537" heatid="4806" lane="3" />
                <RESULT eventid="4429" points="328" swimtime="00:00:32.03" resultid="5568" heatid="4856" lane="3" />
                <RESULT eventid="4431" points="314" swimtime="00:00:32.52" resultid="5574" heatid="4866" lane="3" />
                <RESULT eventid="5807" points="297" swimtime="00:00:37.36" resultid="10286" heatid="6040" lane="7" />
                <RESULT eventid="10332" points="392" swimtime="00:00:27.54" resultid="10506" heatid="10356" lane="1" entrytime="00:00:30.56" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Aparecida Lourenço Alves" birthdate="2013-11-06" gender="F" nation="BRA" license="387374" swrid="5588530" athleteid="3975" externalid="387374" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="151" swimtime="00:00:45.72" resultid="3976" heatid="4664" lane="5" />
                <RESULT eventid="1077" points="198" swimtime="00:00:43.25" resultid="3977" heatid="4715" lane="3" entrytime="00:00:45.39" entrycourse="SCM" />
                <RESULT eventid="1189" status="DNS" swimtime="00:00:00.00" resultid="3978" heatid="4928" lane="3" entrytime="00:01:21.94" entrycourse="SCM" />
                <RESULT eventid="1314" points="238" swimtime="00:00:36.97" resultid="3979" heatid="5088" lane="2" entrytime="00:00:36.74" entrycourse="SCM" />
                <RESULT eventid="1301" points="178" swimtime="00:00:50.35" resultid="3980" heatid="5040" lane="6" entrytime="00:00:57.43" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Luiza Rocha Batista" birthdate="2013-11-24" gender="F" nation="BRA" license="387379" swrid="5588784" athleteid="4002" externalid="387379" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="137" swimtime="00:00:47.24" resultid="4003" heatid="4667" lane="6" entrytime="00:00:46.94" entrycourse="SCM" />
                <RESULT eventid="1077" points="196" swimtime="00:00:43.40" resultid="4004" heatid="4715" lane="2" entrytime="00:00:46.50" entrycourse="SCM" />
                <RESULT eventid="1153" points="129" swimtime="00:01:46.80" resultid="4005" heatid="4900" lane="4" entrytime="00:02:05.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="247" swimtime="00:01:20.00" resultid="4006" heatid="4929" lane="5" entrytime="00:01:19.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="252" swimtime="00:00:36.26" resultid="4007" heatid="5086" lane="7" entrytime="00:00:37.20" entrycourse="SCM" />
                <RESULT eventid="1301" points="95" swimtime="00:01:02.07" resultid="4008" heatid="5032" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Diego" lastname="Brasil Caropreso" birthdate="2009-10-29" gender="M" nation="BRA" license="399502" swrid="5653287" athleteid="4173" externalid="399502" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="355" swimtime="00:00:30.69" resultid="4174" heatid="4779" lane="5" entrytime="00:00:32.28" entrycourse="SCM" />
                <RESULT eventid="1105" points="254" swimtime="00:00:34.89" resultid="4175" heatid="4832" lane="4" />
                <RESULT eventid="1227" points="395" swimtime="00:02:15.38" resultid="4176" heatid="4967" lane="1" entrytime="00:02:14.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.01" />
                    <SPLIT distance="100" swimtime="00:01:01.36" />
                    <SPLIT distance="150" swimtime="00:01:37.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="440" swimtime="00:00:58.95" resultid="4177" heatid="5009" lane="1" entrytime="00:01:01.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="324" swimtime="00:00:36.30" resultid="4179" heatid="5140" lane="1" />
                <RESULT eventid="10332" points="410" swimtime="00:00:27.13" resultid="10536" heatid="10358" lane="4" entrytime="00:00:27.70" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otto" lastname="Hedeke" birthdate="2011-03-24" gender="M" nation="BRA" license="372643" swrid="5588738" athleteid="3913" externalid="372643" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="213" swimtime="00:00:36.40" resultid="3914" heatid="4770" lane="2" />
                <RESULT eventid="1105" points="181" swimtime="00:00:39.07" resultid="3915" heatid="4824" lane="2" />
                <RESULT eventid="1227" points="355" swimtime="00:02:20.26" resultid="3916" heatid="4963" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                    <SPLIT distance="100" swimtime="00:01:08.39" />
                    <SPLIT distance="150" swimtime="00:01:44.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="316" swimtime="00:01:05.83" resultid="3917" heatid="4997" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="227" swimtime="00:00:40.87" resultid="3919" heatid="5140" lane="7" />
                <RESULT eventid="10332" points="291" swimtime="00:00:30.39" resultid="10513" heatid="10351" lane="1" entrytime="00:00:35.55" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabrizio" lastname="Bulla Lanaro" birthdate="2009-08-28" gender="M" nation="BRA" license="344303" swrid="5559846" athleteid="3826" externalid="344303" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="495" swimtime="00:00:27.49" resultid="3827" heatid="4781" lane="5" entrytime="00:00:27.61" entrycourse="SCM" />
                <RESULT eventid="1105" points="412" swimtime="00:00:29.70" resultid="3828" heatid="4825" lane="1" />
                <RESULT eventid="1249" points="361" swimtime="00:01:07.82" resultid="3829" heatid="4983" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1237" points="495" swimtime="00:01:00.37" resultid="3830" heatid="4974" lane="2" entrytime="00:01:02.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="499" swimtime="00:00:31.44" resultid="3832" heatid="5137" lane="3" />
                <RESULT eventid="4423" points="497" swimtime="00:00:27.44" resultid="5547" heatid="4800" lane="1" />
                <RESULT eventid="4425" points="515" swimtime="00:00:27.13" resultid="5553" heatid="4808" lane="1" />
                <RESULT eventid="4429" points="396" swimtime="00:00:30.09" resultid="5587" heatid="4860" lane="3" />
                <RESULT eventid="4431" points="356" swimtime="00:00:31.18" resultid="5602" heatid="4868" lane="3" />
                <RESULT eventid="5807" points="494" swimtime="00:00:31.55" resultid="10296" heatid="6044" lane="5" />
                <RESULT eventid="10332" points="458" swimtime="00:00:26.14" resultid="10502" heatid="10358" lane="7" entrytime="00:00:27.26" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Gelenski Pelaio" birthdate="2005-10-10" gender="M" nation="BRA" license="281473" swrid="5600173" athleteid="3900" externalid="281473" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="583" swimtime="00:00:26.03" resultid="3901" heatid="4781" lane="3" entrytime="00:00:25.91" entrycourse="SCM" />
                <RESULT eventid="4423" points="532" swimtime="00:00:26.84" resultid="5557" heatid="4802" lane="1" />
                <RESULT eventid="4425" points="501" swimtime="00:00:27.38" resultid="5563" heatid="4809" lane="1" />
                <RESULT eventid="10332" points="567" swimtime="00:00:24.35" resultid="10511" heatid="10360" lane="3" entrytime="00:00:24.33" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Victoria De Medeiros" birthdate="2014-08-14" gender="F" nation="BRA" license="403782" swrid="5684611" athleteid="4152" externalid="403782" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="98" swimtime="00:00:52.85" resultid="4153" heatid="4648" lane="4" entrytime="00:00:56.69" entrycourse="SCM" />
                <RESULT eventid="1074" points="86" swimtime="00:00:57.18" resultid="4154" heatid="4697" lane="2" entrytime="00:01:06.21" entrycourse="SCM" />
                <RESULT comment="SW 10.5 - Ao virar, não fez contato com a borda da piscina." eventid="1129" status="DSQ" swimtime="00:02:00.06" resultid="4155" heatid="4881" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="96" swimtime="00:01:57.96" resultid="4156" heatid="4900" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="152" swimtime="00:00:53.10" resultid="4157" heatid="5024" lane="7" entrytime="00:00:58.00" entrycourse="SCM" />
                <RESULT eventid="1311" points="190" swimtime="00:00:39.84" resultid="4158" heatid="5072" lane="3" entrytime="00:00:44.91" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Luiz Cruz" birthdate="2012-10-13" gender="M" nation="BRA" license="393209" swrid="5616447" athleteid="4044" externalid="393209" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="174" swimtime="00:00:38.95" resultid="4045" heatid="4775" lane="5" entrytime="00:00:42.28" entrycourse="SCM" />
                <RESULT eventid="1105" points="102" swimtime="00:00:47.28" resultid="4046" heatid="4824" lane="3" />
                <RESULT eventid="1237" points="113" swimtime="00:01:38.77" resultid="4047" heatid="4970" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="180" swimtime="00:01:19.31" resultid="4048" heatid="4999" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="141" swimtime="00:00:47.88" resultid="4050" heatid="5148" lane="7" entrytime="00:00:49.41" entrycourse="SCM" />
                <RESULT eventid="10332" points="199" swimtime="00:00:34.48" resultid="10525" heatid="10350" lane="8" entrytime="00:00:37.89" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mathias" lastname="Lopes Batista" birthdate="2012-08-22" gender="M" nation="BRA" license="399740" swrid="5652889" athleteid="4085" externalid="399740" level="CLBO">
              <RESULTS>
                <RESULT comment="SW 8.3 - Movimento de pernada de peito.&#10;&#10;&#10;&#10;&#10;&#10;&#10;" eventid="1092" status="DSQ" swimtime="00:00:48.06" resultid="4086" heatid="4769" lane="5" />
                <RESULT eventid="1105" points="165" swimtime="00:00:40.27" resultid="4087" heatid="4836" lane="5" entrytime="00:00:40.85" entrycourse="SCM" />
                <RESULT eventid="1249" points="155" swimtime="00:01:29.93" resultid="4088" heatid="4984" lane="2" entrytime="00:01:39.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="168" swimtime="00:01:21.19" resultid="4089" heatid="5004" lane="1" entrytime="00:01:21.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" status="DNS" swimtime="00:00:00.00" resultid="4091" heatid="5146" lane="2" />
                <RESULT eventid="10332" status="DNS" swimtime="00:00:00.00" resultid="10528" heatid="10351" lane="4" entrytime="00:00:35.30" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Vieira Coelho" birthdate="2014-09-28" gender="F" nation="BRA" license="406951" swrid="5717301" athleteid="4207" externalid="406951" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="124" swimtime="00:00:48.80" resultid="4208" heatid="4650" lane="3" entrytime="00:00:46.69" entrycourse="SCM" />
                <RESULT eventid="1074" points="162" swimtime="00:00:46.25" resultid="4209" heatid="4696" lane="3" />
                <RESULT eventid="1129" points="174" swimtime="00:01:51.66" resultid="4210" heatid="4879" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="154" swimtime="00:01:42.36" resultid="4211" heatid="4911" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" status="DNS" swimtime="00:00:00.00" resultid="4212" heatid="5025" lane="6" entrytime="00:00:52.39" entrycourse="SCM" />
                <RESULT eventid="1311" status="DNS" swimtime="00:00:00.00" resultid="4213" heatid="5072" lane="4" entrytime="00:00:45.77" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Fachini Kovalski" birthdate="2012-05-15" gender="M" nation="BRA" license="403404" swrid="5676297" athleteid="4146" externalid="403404" level="CLBO">
              <RESULTS>
                <RESULT comment="SW 8.3 - Movimento alternado das pernas ou pés." eventid="1092" status="DSQ" swimtime="00:00:54.06" resultid="4147" heatid="4766" lane="2" />
                <RESULT eventid="1105" points="128" swimtime="00:00:43.87" resultid="4148" heatid="4835" lane="3" entrytime="00:00:44.58" entrycourse="SCM" />
                <RESULT eventid="1273" points="127" swimtime="00:01:28.98" resultid="4149" heatid="5002" lane="3" entrytime="00:01:32.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="119" swimtime="00:00:50.68" resultid="4151" heatid="5148" lane="5" entrytime="00:01:01.33" entrycourse="SCM" />
                <RESULT eventid="10332" points="141" swimtime="00:00:38.72" resultid="10535" heatid="10349" lane="2" entrytime="00:00:41.79" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="De Castro Paiva Maciel" birthdate="2008-04-10" gender="M" nation="BRA" license="378333" swrid="5622275" athleteid="3814" externalid="378333" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="493" swimtime="00:00:27.53" resultid="3815" heatid="4780" lane="3" entrytime="00:00:28.95" entrycourse="SCM" />
                <RESULT eventid="1105" points="344" swimtime="00:00:31.54" resultid="3816" heatid="4833" lane="1" />
                <RESULT eventid="1227" points="469" swimtime="00:02:07.86" resultid="3817" heatid="4965" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.38" />
                    <SPLIT distance="100" swimtime="00:01:00.12" />
                    <SPLIT distance="150" swimtime="00:01:34.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="468" swimtime="00:00:57.73" resultid="3818" heatid="5010" lane="5" entrytime="00:00:59.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="292" swimtime="00:00:37.59" resultid="3820" heatid="5146" lane="3" />
                <RESULT eventid="4423" points="505" swimtime="00:00:27.30" resultid="5560" heatid="4802" lane="4" />
                <RESULT eventid="4425" points="454" swimtime="00:00:28.29" resultid="5565" heatid="4809" lane="2" />
                <RESULT eventid="4429" points="348" swimtime="00:00:31.41" resultid="5594" heatid="4862" lane="4" />
                <RESULT eventid="10332" points="468" swimtime="00:00:25.96" resultid="10501" heatid="10359" lane="7" entrytime="00:00:26.82" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucca" lastname="Maceno Araujo" birthdate="2010-09-29" gender="M" nation="BRA" license="367056" swrid="5588788" athleteid="3874" externalid="367056" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="3875" heatid="4779" lane="3" entrytime="00:00:31.01" entrycourse="SCM" />
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="3876" heatid="4829" lane="3" />
                <RESULT eventid="1237" points="351" swimtime="00:01:07.68" resultid="3877" heatid="4974" lane="1" entrytime="00:01:10.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="361" swimtime="00:01:02.97" resultid="3878" heatid="5008" lane="3" entrytime="00:01:02.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="212" swimtime="00:00:41.79" resultid="3880" heatid="5142" lane="2" />
                <RESULT eventid="10332" points="385" swimtime="00:00:27.71" resultid="10507" heatid="10357" lane="6" entrytime="00:00:29.25" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="Soul Santos" birthdate="2016-05-11" gender="M" nation="BRA" license="415247" swrid="5755343" athleteid="4221" externalid="415247" level="CLBO">
              <RESULTS>
                <RESULT eventid="1201" points="51" swimtime="00:00:59.24" resultid="4222" heatid="4940" lane="4" />
                <RESULT eventid="1225" points="32" swimtime="00:01:18.40" resultid="4223" heatid="4960" lane="4" />
                <RESULT eventid="1261" points="75" swimtime="00:00:47.76" resultid="4224" heatid="4990" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Julia Rocha" birthdate="2014-02-10" gender="F" nation="BRA" license="397158" swrid="5641767" athleteid="4057" externalid="397158" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="263" swimtime="00:00:38.04" resultid="4058" heatid="4649" lane="4" entrytime="00:00:53.29" entrycourse="SCM" />
                <RESULT eventid="1074" points="224" swimtime="00:00:41.55" resultid="4059" heatid="4702" lane="3" entrytime="00:00:42.50" entrycourse="SCM" />
                <RESULT eventid="1165" points="230" swimtime="00:01:29.54" resultid="4060" heatid="4908" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="217" swimtime="00:01:29.83" resultid="4061" heatid="4900" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="243" swimtime="00:00:45.41" resultid="4062" heatid="5023" lane="2" entrytime="00:01:01.29" entrycourse="SCM" />
                <RESULT eventid="1311" points="312" swimtime="00:00:33.78" resultid="4063" heatid="5076" lane="2" entrytime="00:00:35.83" entrycourse="SCM" />
                <RESULT eventid="4409" points="273" swimtime="00:00:37.58" resultid="5372" heatid="4656" lane="2" />
                <RESULT eventid="4415" points="231" swimtime="00:00:41.13" resultid="5403" heatid="4707" lane="2" />
                <RESULT eventid="4433" points="257" swimtime="00:00:44.62" resultid="10087" heatid="6064" lane="3" />
                <RESULT eventid="4439" points="318" swimtime="00:00:33.59" resultid="10180" heatid="6050" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lis" lastname="Cristini Harmatiuk" birthdate="2014-07-19" gender="F" nation="BRA" license="396830" swrid="5641759" athleteid="4166" externalid="396830" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="166" swimtime="00:00:44.30" resultid="4167" heatid="4649" lane="2" entrytime="00:00:53.30" entrycourse="SCM" />
                <RESULT eventid="1074" points="186" swimtime="00:00:44.16" resultid="4168" heatid="4702" lane="2" entrytime="00:00:44.65" entrycourse="SCM" />
                <RESULT eventid="1129" points="198" swimtime="00:01:46.82" resultid="4169" heatid="4883" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="171" swimtime="00:01:38.71" resultid="4170" heatid="4905" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" status="DNS" swimtime="00:00:00.00" resultid="4171" heatid="5025" lane="2" entrytime="00:00:50.04" entrycourse="SCM" />
                <RESULT eventid="1311" status="DNS" swimtime="00:00:00.00" resultid="4172" heatid="5075" lane="7" entrytime="00:00:41.73" entrycourse="SCM" />
                <RESULT eventid="4409" points="159" swimtime="00:00:44.98" resultid="5373" heatid="4656" lane="5" />
                <RESULT eventid="4415" points="197" swimtime="00:00:43.34" resultid="5406" heatid="4707" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Marcos Morais" birthdate="2010-01-30" gender="M" nation="BRA" license="416736" swrid="5757093" athleteid="4244" externalid="416736" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="279" swimtime="00:00:33.28" resultid="4245" heatid="4770" lane="3" />
                <RESULT eventid="1105" points="244" swimtime="00:00:35.38" resultid="4246" heatid="4826" lane="2" />
                <RESULT eventid="1213" points="328" swimtime="00:01:20.08" resultid="4247" heatid="4950" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="304" swimtime="00:01:06.64" resultid="4248" heatid="4997" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="320" swimtime="00:00:36.45" resultid="4250" heatid="5142" lane="8" />
                <RESULT eventid="4429" points="253" swimtime="00:00:34.93" resultid="5581" heatid="4858" lane="6" />
                <RESULT eventid="5807" points="341" swimtime="00:00:35.69" resultid="10291" heatid="6042" lane="7" />
                <RESULT eventid="10332" points="330" swimtime="00:00:29.15" resultid="10541" heatid="10347" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Prestes Alves Pinto" birthdate="2012-01-19" gender="F" nation="BRA" license="377324" swrid="5588867" athleteid="3947" externalid="377324" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="276" swimtime="00:00:37.42" resultid="3948" heatid="4662" lane="6" />
                <RESULT eventid="1077" points="291" swimtime="00:00:38.08" resultid="3949" heatid="4720" lane="3" entrytime="00:00:37.14" entrycourse="SCM" />
                <RESULT eventid="1119" points="301" swimtime="00:02:57.43" resultid="3950" heatid="4876" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                    <SPLIT distance="100" swimtime="00:01:25.19" />
                    <SPLIT distance="150" swimtime="00:02:11.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="371" swimtime="00:02:33.40" resultid="3951" heatid="4895" lane="1" entrytime="00:02:40.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.78" />
                    <SPLIT distance="100" swimtime="00:01:14.00" />
                    <SPLIT distance="150" swimtime="00:01:54.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="398" swimtime="00:00:31.16" resultid="3952" heatid="5090" lane="2" entrytime="00:00:33.87" entrycourse="SCM" />
                <RESULT eventid="1301" points="219" swimtime="00:00:47.00" resultid="3953" heatid="5032" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Zanotto Souza" birthdate="2015-07-01" gender="M" nation="BRA" license="415249" swrid="5755347" athleteid="4225" externalid="415249" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="49" swimtime="00:00:59.19" resultid="4226" heatid="4750" lane="5" />
                <RESULT eventid="1102" status="DSQ" swimtime="00:00:54.02" resultid="4227" heatid="4811" lane="4" />
                <RESULT eventid="1273" points="85" swimtime="00:01:41.89" resultid="4228" heatid="5000" lane="2" />
                <RESULT eventid="1326" points="60" swimtime="00:01:03.70" resultid="4230" heatid="5127" lane="8" />
                <RESULT eventid="10329" points="106" swimtime="00:00:42.55" resultid="10539" heatid="10341" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Breno" lastname="Borges Piekarzievicz" birthdate="2011-11-11" gender="M" nation="BRA" license="403144" swrid="5676295" athleteid="4132" externalid="403144" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="4133" heatid="4767" lane="4" />
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="4134" heatid="4834" lane="2" />
                <RESULT eventid="1213" status="DNS" swimtime="00:00:00.00" resultid="4135" heatid="4950" lane="1" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="4136" heatid="5001" lane="6" />
                <RESULT eventid="1329" points="145" swimtime="00:00:47.43" resultid="4138" heatid="5139" lane="2" />
                <RESULT eventid="10332" points="183" swimtime="00:00:35.49" resultid="10534" heatid="10349" lane="3" entrytime="00:00:40.55" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tais" lastname="Feltrin Martins" birthdate="2013-01-17" gender="F" nation="BRA" license="406840" swrid="5717262" athleteid="4180" externalid="406840" level="CLBO">
              <RESULTS>
                <RESULT comment="SW 8.5 - Totalmente submerso durante o nado." eventid="1064" status="DSQ" swimtime="00:01:16.01" resultid="4181" heatid="4660" lane="4" />
                <RESULT eventid="1077" points="87" swimtime="00:00:56.77" resultid="4182" heatid="4714" lane="4" entrytime="00:00:57.24" entrycourse="SCM" />
                <RESULT eventid="1165" points="85" swimtime="00:02:04.61" resultid="4183" heatid="4912" lane="6" entrytime="00:02:10.57" entrycourse="SCM" />
                <RESULT eventid="1314" points="114" swimtime="00:00:47.22" resultid="4184" heatid="5085" lane="3" entrytime="00:00:46.58" entrycourse="SCM" />
                <RESULT eventid="1301" points="74" swimtime="00:01:07.38" resultid="4185" heatid="5038" lane="3" entrytime="00:01:07.54" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Zanotto De Souza" birthdate="2013-08-24" gender="M" nation="BRA" license="388361" swrid="5588974" athleteid="4016" externalid="388361" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="217" swimtime="00:00:36.17" resultid="4017" heatid="4772" lane="1" />
                <RESULT eventid="1105" points="165" swimtime="00:00:40.29" resultid="4018" heatid="4837" lane="6" entrytime="00:00:39.69" entrycourse="SCM" />
                <RESULT eventid="1237" points="156" swimtime="00:01:28.61" resultid="4019" heatid="4970" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="224" swimtime="00:01:13.78" resultid="4020" heatid="5006" lane="5" entrytime="00:01:12.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="149" swimtime="00:00:47.02" resultid="4022" heatid="5150" lane="6" entrytime="00:00:49.33" entrycourse="SCM" />
                <RESULT eventid="4425" points="186" swimtime="00:00:38.08" resultid="5478" heatid="4804" lane="3" />
                <RESULT eventid="4423" points="220" swimtime="00:00:36.01" resultid="5484" heatid="4792" lane="4" />
                <RESULT eventid="4429" points="195" swimtime="00:00:38.10" resultid="5516" heatid="4852" lane="6" />
                <RESULT eventid="4431" points="151" swimtime="00:00:41.43" resultid="5517" heatid="4864" lane="1" />
                <RESULT eventid="10332" points="256" swimtime="00:00:31.72" resultid="10521" heatid="10354" lane="1" entrytime="00:00:31.95" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Augusto Vaz" birthdate="2011-06-25" gender="M" nation="BRA" license="401737" swrid="5661339" athleteid="4113" externalid="401737" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="429" swimtime="00:00:28.82" resultid="4114" heatid="4776" lane="3" entrytime="00:00:37.52" entrycourse="SCM" />
                <RESULT eventid="1105" points="286" swimtime="00:00:33.55" resultid="4115" heatid="4832" lane="5" />
                <RESULT eventid="1237" points="397" swimtime="00:01:05.00" resultid="4116" heatid="4971" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="392" swimtime="00:01:01.24" resultid="4117" heatid="4996" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="217" swimtime="00:00:41.50" resultid="4119" heatid="5140" lane="5" />
                <RESULT eventid="4423" points="421" swimtime="00:00:29.00" resultid="5529" heatid="4796" lane="1" />
                <RESULT eventid="4425" points="354" swimtime="00:00:30.74" resultid="5535" heatid="4806" lane="1" />
                <RESULT eventid="4429" points="322" swimtime="00:00:32.23" resultid="5569" heatid="4856" lane="4" />
                <RESULT eventid="10332" points="385" swimtime="00:00:27.69" resultid="10531" heatid="10354" lane="8" entrytime="00:00:32.38" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabio" lastname="C Burak" birthdate="2009-08-29" gender="M" nation="BRA" license="343297" swrid="5600126" athleteid="4037" externalid="343297" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="456" swimtime="00:00:28.25" resultid="4038" heatid="4770" lane="4" />
                <RESULT eventid="1105" points="432" swimtime="00:00:29.23" resultid="4039" heatid="4828" lane="4" />
                <RESULT eventid="1249" points="479" swimtime="00:01:01.75" resultid="4040" heatid="4986" lane="4" entrytime="00:01:04.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1237" status="DNS" swimtime="00:00:00.00" resultid="4041" heatid="4971" lane="2" />
                <RESULT eventid="1329" points="465" swimtime="00:00:32.19" resultid="4043" heatid="5155" lane="5" entrytime="00:00:33.15" entrycourse="SCM" />
                <RESULT eventid="4423" points="487" swimtime="00:00:27.63" resultid="5550" heatid="4800" lane="4" />
                <RESULT eventid="4425" points="405" swimtime="00:00:29.38" resultid="5555" heatid="4808" lane="3" />
                <RESULT eventid="4429" points="433" swimtime="00:00:29.22" resultid="5585" heatid="4860" lane="1" />
                <RESULT eventid="4431" points="410" swimtime="00:00:29.75" resultid="5600" heatid="4868" lane="1" />
                <RESULT eventid="5807" points="472" swimtime="00:00:32.04" resultid="10297" heatid="6044" lane="6" />
                <RESULT eventid="10332" points="475" swimtime="00:00:25.82" resultid="10524" heatid="10358" lane="1" entrytime="00:00:27.91" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Analyce" lastname="Nunes Porto Luz" birthdate="2006-10-29" gender="F" nation="BRA" license="369322" swrid="5600226" athleteid="3811" externalid="369322" level="CLBO">
              <RESULTS>
                <RESULT eventid="1314" points="519" swimtime="00:00:28.53" resultid="3813" heatid="5084" lane="3" />
                <RESULT eventid="1064" points="463" swimtime="00:00:31.51" resultid="5255" heatid="4657" lane="6" />
                <RESULT eventid="1077" points="383" swimtime="00:00:34.75" resultid="5325" heatid="4714" lane="1" />
                <RESULT eventid="4411" points="450" swimtime="00:00:31.80" resultid="5344" heatid="4688" lane="1" />
                <RESULT eventid="4413" points="406" swimtime="00:00:32.92" resultid="5350" heatid="4695" lane="1" />
                <RESULT eventid="4417" points="393" swimtime="00:00:34.45" resultid="5454" heatid="4739" lane="1" />
                <RESULT eventid="4419" points="395" swimtime="00:00:34.41" resultid="5460" heatid="4746" lane="1" />
                <RESULT eventid="5804" points="511" swimtime="00:00:28.68" resultid="10218" heatid="6062" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Rodrigues Bortoluzzi" birthdate="2013-10-07" gender="M" nation="BRA" license="387375" swrid="5652897" athleteid="3981" externalid="387375" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="136" swimtime="00:00:42.27" resultid="3982" heatid="4774" lane="1" />
                <RESULT eventid="1105" points="141" swimtime="00:00:42.47" resultid="3983" heatid="4835" lane="6" entrytime="00:00:46.67" entrycourse="SCM" />
                <RESULT eventid="1203" points="157" swimtime="00:03:15.54" resultid="3984" heatid="4942" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.00" />
                    <SPLIT distance="100" swimtime="00:01:35.12" />
                    <SPLIT distance="150" swimtime="00:02:26.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="145" swimtime="00:01:31.85" resultid="3985" heatid="4984" lane="1" entrytime="00:01:50.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="100" swimtime="00:00:53.63" resultid="3987" heatid="5148" lane="1" entrytime="00:01:03.02" entrycourse="SCM" />
                <RESULT eventid="10332" points="182" swimtime="00:00:35.51" resultid="10517" heatid="10350" lane="6" entrytime="00:00:36.99" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lauren" lastname="Kurecki" birthdate="2014-03-06" gender="F" nation="BRA" license="377314" swrid="5602549" athleteid="3927" externalid="377314" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="250" swimtime="00:00:38.70" resultid="3928" heatid="4651" lane="2" entrytime="00:00:41.26" entrycourse="SCM" />
                <RESULT eventid="1074" points="195" swimtime="00:00:43.49" resultid="3929" heatid="4697" lane="6" />
                <RESULT eventid="1129" points="261" swimtime="00:01:37.50" resultid="3930" heatid="4884" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="281" swimtime="00:01:16.70" resultid="3931" heatid="4930" lane="2" entrytime="00:01:13.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="262" swimtime="00:00:44.32" resultid="3932" heatid="5025" lane="3" entrytime="00:00:43.37" entrycourse="SCM" />
                <RESULT eventid="1311" points="300" swimtime="00:00:34.23" resultid="3933" heatid="5076" lane="3" entrytime="00:00:33.10" entrycourse="SCM" />
                <RESULT eventid="4409" points="242" swimtime="00:00:39.10" resultid="5370" heatid="4656" lane="3" />
                <RESULT eventid="4415" points="213" swimtime="00:00:42.22" resultid="5404" heatid="4707" lane="3" />
                <RESULT eventid="4433" points="285" swimtime="00:00:43.06" resultid="10085" heatid="6064" lane="1" />
                <RESULT eventid="4439" points="325" swimtime="00:00:33.34" resultid="10181" heatid="6050" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Victor Dallastra" birthdate="2010-08-21" gender="M" nation="BRA" license="408024" swrid="5723028" athleteid="4214" externalid="408024" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="334" swimtime="00:00:31.32" resultid="4215" heatid="4762" lane="2" />
                <RESULT eventid="1105" points="195" swimtime="00:00:38.07" resultid="4216" heatid="4832" lane="1" />
                <RESULT eventid="1227" points="422" swimtime="00:02:12.41" resultid="4217" heatid="4962" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.02" />
                    <SPLIT distance="100" swimtime="00:01:01.21" />
                    <SPLIT distance="150" swimtime="00:01:36.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="390" swimtime="00:01:01.34" resultid="4218" heatid="5000" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="278" swimtime="00:00:38.19" resultid="4220" heatid="5146" lane="6" />
                <RESULT eventid="4423" points="313" swimtime="00:00:32.00" resultid="5542" heatid="4798" lane="5" />
                <RESULT eventid="10332" points="384" swimtime="00:00:27.72" resultid="10538" heatid="10348" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Bulla Lanaro" birthdate="2009-08-28" gender="F" nation="BRA" license="344301" swrid="5569976" athleteid="3801" externalid="344301" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="556" swimtime="00:00:29.64" resultid="3802" heatid="4671" lane="3" entrytime="00:00:31.21" entrycourse="SCM" />
                <RESULT eventid="1077" points="496" swimtime="00:00:31.88" resultid="3803" heatid="4713" lane="4" />
                <RESULT eventid="1165" points="477" swimtime="00:01:10.22" resultid="3804" heatid="4907" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="566" swimtime="00:01:05.32" resultid="3805" heatid="4901" lane="3" entrytime="00:01:05.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="585" swimtime="00:01:00.06" resultid="3806" heatid="4933" lane="3" entrytime="00:01:01.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="559" swimtime="00:00:27.83" resultid="3807" heatid="5097" lane="3" entrytime="00:00:27.94" entrycourse="SCM" />
                <RESULT eventid="4411" points="531" swimtime="00:00:30.10" resultid="5335" heatid="4686" lane="1" />
                <RESULT eventid="4413" points="508" swimtime="00:00:30.54" resultid="5341" heatid="4694" lane="1" />
                <RESULT eventid="4417" points="448" swimtime="00:00:32.98" resultid="5445" heatid="4737" lane="1" />
                <RESULT eventid="4419" points="490" swimtime="00:00:32.01" resultid="5451" heatid="4745" lane="1" />
                <RESULT eventid="5804" points="567" swimtime="00:00:27.69" resultid="10212" heatid="6060" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lais" lastname="Manika Broto" birthdate="2013-03-27" gender="F" nation="BRA" license="378054" swrid="5588795" athleteid="3954" externalid="378054" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="331" swimtime="00:00:35.23" resultid="3955" heatid="4670" lane="5" entrytime="00:00:36.63" entrycourse="SCM" />
                <RESULT eventid="1077" points="263" swimtime="00:00:39.37" resultid="3956" heatid="4713" lane="5" />
                <RESULT eventid="1153" points="257" swimtime="00:01:24.99" resultid="3957" heatid="4899" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="389" swimtime="00:01:08.81" resultid="3958" heatid="4931" lane="3" entrytime="00:01:09.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="389" swimtime="00:00:31.40" resultid="3959" heatid="5089" lane="3" entrytime="00:00:35.10" entrycourse="SCM" />
                <RESULT eventid="1301" points="228" swimtime="00:00:46.40" resultid="3960" heatid="5034" lane="3" />
                <RESULT eventid="4413" points="307" swimtime="00:00:36.12" resultid="5376" heatid="4690" lane="2" />
                <RESULT eventid="4411" points="332" swimtime="00:00:35.20" resultid="5382" heatid="4678" lane="2" />
                <RESULT eventid="4417" points="280" swimtime="00:00:38.57" resultid="5412" heatid="4729" lane="5" />
                <RESULT eventid="5804" points="402" swimtime="00:00:31.05" resultid="10187" heatid="6052" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Marques" birthdate="2007-06-29" gender="M" nation="BRA" license="367257" swrid="5600213" athleteid="4200" externalid="367257" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="293" swimtime="00:00:32.72" resultid="4201" heatid="4762" lane="4" />
                <RESULT eventid="1105" points="204" swimtime="00:00:37.55" resultid="4202" heatid="4830" lane="1" />
                <RESULT eventid="1227" points="321" swimtime="00:02:25.02" resultid="4203" heatid="4963" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                    <SPLIT distance="100" swimtime="00:01:09.04" />
                    <SPLIT distance="150" swimtime="00:01:47.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="317" swimtime="00:01:05.73" resultid="4204" heatid="5008" lane="2" entrytime="00:01:03.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="185" swimtime="00:00:43.71" resultid="4206" heatid="5143" lane="7" />
                <RESULT eventid="10332" points="339" swimtime="00:00:28.90" resultid="10537" heatid="10347" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Nogueira Silva" birthdate="2011-08-13" gender="M" nation="BRA" license="367150" swrid="5588832" athleteid="3888" externalid="367150" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="244" swimtime="00:00:34.77" resultid="3889" heatid="4772" lane="2" />
                <RESULT eventid="1105" points="189" swimtime="00:00:38.48" resultid="3890" heatid="4831" lane="6" />
                <RESULT eventid="1227" points="353" swimtime="00:02:20.53" resultid="3891" heatid="4965" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:01:07.11" />
                    <SPLIT distance="150" swimtime="00:01:44.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="308" swimtime="00:01:06.35" resultid="3892" heatid="4996" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="284" swimtime="00:00:37.92" resultid="3894" heatid="5139" lane="7" />
                <RESULT eventid="5807" points="285" swimtime="00:00:37.89" resultid="10279" heatid="6040" lane="2" />
                <RESULT eventid="10332" points="328" swimtime="00:00:29.22" resultid="10509" heatid="10356" lane="2" entrytime="00:00:30.27" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Guilherme Ieger" birthdate="2009-02-20" gender="M" nation="BRA" license="356888" swrid="5600180" athleteid="3853" externalid="356888" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="370" swimtime="00:00:30.27" resultid="3854" heatid="4773" lane="1" />
                <RESULT eventid="1105" points="289" swimtime="00:00:33.43" resultid="3855" heatid="4831" lane="3" />
                <RESULT eventid="1213" points="412" swimtime="00:01:14.26" resultid="3856" heatid="4954" lane="2" entrytime="00:01:15.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="449" swimtime="00:00:58.54" resultid="3857" heatid="5010" lane="1" entrytime="00:01:00.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="425" swimtime="00:00:33.16" resultid="3859" heatid="5155" lane="6" entrytime="00:00:35.32" entrycourse="SCM" />
                <RESULT eventid="5807" points="422" swimtime="00:00:33.24" resultid="10293" heatid="6044" lane="2" />
                <RESULT eventid="10332" points="447" swimtime="00:00:26.35" resultid="10505" heatid="10359" lane="1" entrytime="00:00:26.62" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mathias" lastname="Bernardo" birthdate="2014-05-17" gender="M" nation="BRA" license="387376" swrid="5652880" athleteid="3988" externalid="387376" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="88" swimtime="00:00:48.85" resultid="3989" heatid="4751" lane="4" />
                <RESULT eventid="1102" points="82" swimtime="00:00:50.82" resultid="3990" heatid="4815" lane="3" entrytime="00:00:49.40" entrycourse="SCM" />
                <RESULT eventid="1249" points="94" swimtime="00:01:46.27" resultid="3991" heatid="4980" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="133" swimtime="00:01:27.64" resultid="3992" heatid="5002" lane="1" entrytime="00:01:39.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="95" swimtime="00:00:54.59" resultid="3994" heatid="5130" lane="8" entrytime="00:00:58.50" entrycourse="SCM" />
                <RESULT eventid="10329" points="154" swimtime="00:00:37.56" resultid="10518" heatid="10343" lane="4" entrytime="00:00:40.10" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Zattar" birthdate="2012-04-19" gender="F" nation="BRA" license="401736" swrid="5661351" athleteid="4106" externalid="401736" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="359" swimtime="00:00:34.29" resultid="4107" heatid="4662" lane="2" />
                <RESULT eventid="1077" points="319" swimtime="00:00:36.92" resultid="4108" heatid="4718" lane="4" entrytime="00:00:40.35" entrycourse="SCM" />
                <RESULT eventid="1119" points="257" swimtime="00:03:07.00" resultid="4109" heatid="4876" lane="6" />
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 5:50), Na volta dos 50m." eventid="1179" status="DSQ" swimtime="00:03:17.97" resultid="4110" heatid="4922" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                    <SPLIT distance="100" swimtime="00:01:32.00" />
                    <SPLIT distance="150" swimtime="00:02:25.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="382" swimtime="00:00:31.60" resultid="4111" heatid="5089" lane="7" entrytime="00:00:36.44" entrycourse="SCM" />
                <RESULT eventid="1301" points="348" swimtime="00:00:40.32" resultid="4112" heatid="5034" lane="1" />
                <RESULT eventid="4411" points="349" swimtime="00:00:34.61" resultid="5390" heatid="4680" lane="4" />
                <RESULT eventid="4417" points="305" swimtime="00:00:37.49" resultid="5422" heatid="4731" lane="6" />
                <RESULT eventid="5801" points="346" swimtime="00:00:40.41" resultid="10098" heatid="6068" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juliana" lastname="Cirilo Da Cunha" birthdate="2013-05-26" gender="F" nation="BRA" license="377316" swrid="5588595" athleteid="3934" externalid="377316" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="258" swimtime="00:00:38.25" resultid="3935" heatid="4663" lane="6" />
                <RESULT eventid="1077" points="236" swimtime="00:00:40.85" resultid="3936" heatid="4709" lane="4" />
                <RESULT eventid="1189" status="DNS" swimtime="00:00:00.00" resultid="3937" heatid="4929" lane="1" entrytime="00:01:19.86" entrycourse="SCM" />
                <RESULT eventid="1314" points="289" swimtime="00:00:34.65" resultid="3938" heatid="5089" lane="6" entrytime="00:00:35.44" entrycourse="SCM" />
                <RESULT eventid="1301" points="198" swimtime="00:00:48.67" resultid="3939" heatid="5041" lane="7" entrytime="00:00:55.86" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Hugo Dos Santos" birthdate="2014-07-25" gender="M" nation="BRA" license="397420" swrid="5641766" athleteid="4071" externalid="397420" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="121" swimtime="00:00:43.92" resultid="4072" heatid="4755" lane="6" entrytime="00:00:49.40" entrycourse="SCM" />
                <RESULT eventid="1102" points="109" swimtime="00:00:46.22" resultid="4073" heatid="4814" lane="3" entrytime="00:00:52.62" entrycourse="SCM" />
                <RESULT eventid="1213" points="124" swimtime="00:01:50.73" resultid="4074" heatid="4951" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="117" swimtime="00:01:38.63" resultid="4075" heatid="4980" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="118" swimtime="00:00:50.82" resultid="4077" heatid="5128" lane="2" entrytime="00:01:02.05" entrycourse="SCM" />
                <RESULT eventid="10329" points="178" swimtime="00:00:35.78" resultid="10526" heatid="10343" lane="2" entrytime="00:00:40.11" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexandre" lastname="Prestes" birthdate="2014-01-16" gender="M" nation="BRA" license="382249" swrid="5602574" athleteid="3968" externalid="382249" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="102" swimtime="00:00:46.41" resultid="3969" heatid="4754" lane="5" entrytime="00:00:54.09" entrycourse="SCM" />
                <RESULT eventid="1102" points="106" swimtime="00:00:46.66" resultid="3970" heatid="4817" lane="6" entrytime="00:00:43.09" entrycourse="SCM" />
                <RESULT eventid="1213" points="151" swimtime="00:01:43.64" resultid="3971" heatid="4947" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="158" swimtime="00:01:22.92" resultid="3972" heatid="5004" lane="6" entrytime="00:01:23.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="159" swimtime="00:00:45.96" resultid="3974" heatid="5131" lane="2" entrytime="00:00:48.48" entrycourse="SCM" />
                <RESULT eventid="4445" points="149" swimtime="00:00:47.02" resultid="10313" heatid="6034" lane="3" />
                <RESULT eventid="10329" points="187" swimtime="00:00:35.22" resultid="10516" heatid="10345" lane="1" entrytime="00:00:36.04" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cleverson" lastname="Cardoso" birthdate="2013-07-20" gender="M" nation="BRA" license="387382" swrid="5588577" athleteid="4009" externalid="387382" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="121" swimtime="00:00:43.90" resultid="4010" heatid="4770" lane="5" />
                <RESULT eventid="1105" points="120" swimtime="00:00:44.73" resultid="4011" heatid="4835" lane="5" entrytime="00:00:46.41" entrycourse="SCM" />
                <RESULT eventid="1263" points="165" swimtime="00:03:38.80" resultid="4012" heatid="4992" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.08" />
                    <SPLIT distance="100" swimtime="00:01:45.34" />
                    <SPLIT distance="150" swimtime="00:02:42.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="184" swimtime="00:01:18.73" resultid="4013" heatid="5003" lane="4" entrytime="00:01:25.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="159" swimtime="00:00:45.96" resultid="4015" heatid="5150" lane="2" entrytime="00:00:51.23" entrycourse="SCM" />
                <RESULT eventid="5807" points="151" swimtime="00:00:46.78" resultid="10272" heatid="6036" lane="7" />
                <RESULT eventid="10332" points="190" swimtime="00:00:35.03" resultid="10520" heatid="10350" lane="1" entrytime="00:00:38.90" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Gabriel Broto" birthdate="2014-09-14" gender="M" nation="BRA" license="402171" swrid="5661345" athleteid="4120" externalid="402171" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="31" swimtime="00:01:08.72" resultid="4121" heatid="4751" lane="3" />
                <RESULT eventid="1102" points="47" swimtime="00:01:01.21" resultid="4122" heatid="4813" lane="5" entrytime="00:01:01.75" entrycourse="SCM" />
                <RESULT eventid="1326" status="DNS" swimtime="00:00:00.00" resultid="4124" heatid="5126" lane="4" />
                <RESULT eventid="10329" status="DNS" swimtime="00:00:00.00" resultid="10532" heatid="10341" lane="5" entrytime="00:00:51.78" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Ryan Rosa" birthdate="2014-01-14" gender="M" nation="BRA" license="400032" swrid="5652898" athleteid="4099" externalid="400032" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="54" swimtime="00:00:57.48" resultid="4100" heatid="4749" lane="3" />
                <RESULT eventid="1102" points="96" swimtime="00:00:48.26" resultid="4101" heatid="4816" lane="6" entrytime="00:00:49.01" entrycourse="SCM" />
                <RESULT eventid="1213" points="114" swimtime="00:01:53.68" resultid="4102" heatid="4946" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="118" swimtime="00:01:31.24" resultid="4103" heatid="5002" lane="4" entrytime="00:01:32.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="100" swimtime="00:00:53.68" resultid="4105" heatid="5130" lane="3" entrytime="00:00:52.86" entrycourse="SCM" />
                <RESULT eventid="10329" points="133" swimtime="00:00:39.43" resultid="10530" heatid="10343" lane="8" entrytime="00:00:39.45" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helloisa" lastname="De Bassani" birthdate="2012-09-23" gender="F" nation="BRA" license="403403" swrid="5676296" athleteid="4139" externalid="403403" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="80" swimtime="00:00:56.42" resultid="4140" heatid="4657" lane="4" />
                <RESULT eventid="1077" points="126" swimtime="00:00:50.27" resultid="4141" heatid="4715" lane="1" entrytime="00:00:50.33" entrycourse="SCM" />
                <RESULT eventid="1129" points="108" swimtime="00:02:10.78" resultid="4142" heatid="4884" lane="4" entrytime="00:02:39.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="157" swimtime="00:01:33.05" resultid="4143" heatid="4927" lane="2" entrytime="00:01:35.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="186" swimtime="00:00:40.12" resultid="4144" heatid="5086" lane="6" entrytime="00:00:41.10" entrycourse="SCM" />
                <RESULT eventid="1301" points="121" swimtime="00:00:57.33" resultid="4145" heatid="5038" lane="7" entrytime="00:00:59.38" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kethelyn" lastname="Ribeiro Rodrigues" birthdate="2009-04-24" gender="F" nation="BRA" license="367052" swrid="5600244" athleteid="3860" externalid="367052" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="277" swimtime="00:00:37.40" resultid="3861" heatid="4658" lane="3" />
                <RESULT eventid="1077" points="270" swimtime="00:00:39.02" resultid="3862" heatid="4720" lane="6" entrytime="00:00:38.51" entrycourse="SCM" />
                <RESULT eventid="1165" points="272" swimtime="00:01:24.69" resultid="3863" heatid="4904" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="389" swimtime="00:01:08.81" resultid="3864" heatid="4932" lane="5" entrytime="00:01:07.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="399" swimtime="00:00:31.13" resultid="3865" heatid="5096" lane="7" entrytime="00:00:30.69" entrycourse="SCM" />
                <RESULT eventid="1301" points="209" swimtime="00:00:47.74" resultid="3866" heatid="5037" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Lopes Rempel" birthdate="2010-09-25" gender="M" nation="BRA" license="399739" swrid="5653294" athleteid="4078" externalid="399739" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="228" swimtime="00:00:35.56" resultid="4079" heatid="4768" lane="6" />
                <RESULT eventid="1105" points="256" swimtime="00:00:34.79" resultid="4080" heatid="4838" lane="4" entrytime="00:00:37.06" entrycourse="SCM" />
                <RESULT eventid="1249" points="254" swimtime="00:01:16.23" resultid="4081" heatid="4985" lane="5" entrytime="00:01:24.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="273" swimtime="00:01:09.06" resultid="4082" heatid="4997" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="171" swimtime="00:00:44.92" resultid="4084" heatid="5143" lane="8" />
                <RESULT eventid="4429" points="266" swimtime="00:00:34.37" resultid="5580" heatid="4858" lane="5" />
                <RESULT eventid="10332" points="291" swimtime="00:00:30.42" resultid="10527" heatid="10354" lane="6" entrytime="00:00:31.96" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Novakoski" birthdate="2009-03-05" gender="F" nation="BRA" license="339136" swrid="5600225" athleteid="3840" externalid="339136" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="419" swimtime="00:00:32.57" resultid="3841" heatid="4665" lane="4" />
                <RESULT eventid="1077" points="296" swimtime="00:00:37.86" resultid="3842" heatid="4708" lane="4" />
                <RESULT eventid="1189" points="494" swimtime="00:01:03.55" resultid="3843" heatid="4932" lane="3" entrytime="00:01:06.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="475" swimtime="00:00:29.38" resultid="3844" heatid="5094" lane="8" entrytime="00:00:30.62" entrycourse="SCM" />
                <RESULT comment="SW 7.1 - Mais de uma pernada de borboleta antes da primeira pernada de peito após o início ou a virada., Após a volta dos 25m." eventid="1301" status="DSQ" swimtime="00:00:44.13" resultid="3845" heatid="5036" lane="4" />
                <RESULT eventid="4411" points="403" swimtime="00:00:32.99" resultid="5338" heatid="4686" lane="4" />
                <RESULT eventid="4417" points="334" swimtime="00:00:36.39" resultid="5450" heatid="4737" lane="6" />
                <RESULT eventid="4423" points="287" swimtime="00:00:36.93" resultid="5703" heatid="4795" lane="5" />
                <RESULT eventid="5804" points="443" swimtime="00:00:30.06" resultid="10211" heatid="6060" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Cavassin Ieger" birthdate="2011-08-31" gender="M" nation="BRA" license="367149" swrid="5588743" athleteid="3881" externalid="367149" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="288" swimtime="00:00:32.90" resultid="3882" heatid="4767" lane="5" />
                <RESULT eventid="1105" points="228" swimtime="00:00:36.14" resultid="3883" heatid="4827" lane="1" />
                <RESULT eventid="1213" points="295" swimtime="00:01:22.97" resultid="3884" heatid="4953" lane="5" entrytime="00:01:26.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="303" swimtime="00:02:58.72" resultid="3885" heatid="4993" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.56" />
                    <SPLIT distance="100" swimtime="00:01:25.71" />
                    <SPLIT distance="150" swimtime="00:02:12.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="287" swimtime="00:00:37.81" resultid="3887" heatid="5154" lane="2" entrytime="00:00:38.96" entrycourse="SCM" />
                <RESULT eventid="5807" points="276" swimtime="00:00:38.29" resultid="10284" heatid="6040" lane="6" />
                <RESULT eventid="10332" points="273" swimtime="00:00:31.07" resultid="10508" heatid="10353" lane="8" entrytime="00:00:33.42" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1115" points="298" swimtime="00:04:28.57" resultid="4259" heatid="4871" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                    <SPLIT distance="100" swimtime="00:01:12.03" />
                    <SPLIT distance="150" swimtime="00:01:43.31" />
                    <SPLIT distance="200" swimtime="00:02:20.20" />
                    <SPLIT distance="250" swimtime="00:02:48.16" />
                    <SPLIT distance="300" swimtime="00:03:25.54" />
                    <SPLIT distance="350" swimtime="00:04:01.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4023" number="1" />
                    <RELAYPOSITION athleteid="3968" number="2" />
                    <RELAYPOSITION athleteid="4016" number="3" />
                    <RELAYPOSITION athleteid="3903" number="4" />
                    <RELAYPOSITION athleteid="3867" number="5" />
                    <RELAYPOSITION athleteid="4244" number="6" />
                    <RELAYPOSITION athleteid="3826" number="7" />
                    <RELAYPOSITION athleteid="3814" number="8" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1339" points="323" swimtime="00:03:58.44" resultid="4260" heatid="5246" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                    <SPLIT distance="100" swimtime="00:01:10.90" />
                    <SPLIT distance="150" swimtime="00:01:42.97" />
                    <SPLIT distance="200" swimtime="00:02:12.23" />
                    <SPLIT distance="250" swimtime="00:02:39.85" />
                    <SPLIT distance="300" swimtime="00:03:07.28" />
                    <SPLIT distance="350" swimtime="00:03:33.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4023" number="1" />
                    <RELAYPOSITION athleteid="3968" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4016" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3903" number="4" reactiontime="0" />
                    <RELAYPOSITION athleteid="3867" number="5" reactiontime="0" />
                    <RELAYPOSITION athleteid="4214" number="6" reactiontime="0" />
                    <RELAYPOSITION athleteid="3826" number="7" reactiontime="0" />
                    <RELAYPOSITION athleteid="3814" number="8" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida." eventid="1087" status="DSQ" swimtime="00:04:53.24" resultid="4257" heatid="4748" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3927" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="3954" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="4106" number="4" status="DSQ" />
                    <RELAYPOSITION athleteid="4159" number="5" status="DSQ" />
                    <RELAYPOSITION athleteid="4186" number="6" status="DSQ" />
                    <RELAYPOSITION athleteid="3801" number="7" status="DSQ" />
                    <RELAYPOSITION athleteid="3811" number="8" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1324" points="378" swimtime="00:04:15.82" resultid="4258" heatid="5123" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="100" swimtime="00:01:06.22" />
                    <SPLIT distance="150" swimtime="00:01:37.08" />
                    <SPLIT distance="200" swimtime="00:02:13.99" />
                    <SPLIT distance="250" swimtime="00:02:48.35" />
                    <SPLIT distance="300" swimtime="00:03:19.52" />
                    <SPLIT distance="350" swimtime="00:03:47.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3927" number="1" />
                    <RELAYPOSITION number="2" />
                    <RELAYPOSITION athleteid="3954" number="3" />
                    <RELAYPOSITION athleteid="4106" number="4" />
                    <RELAYPOSITION athleteid="4159" number="5" />
                    <RELAYPOSITION athleteid="4186" number="6" />
                    <RELAYPOSITION athleteid="3801" number="7" />
                    <RELAYPOSITION athleteid="3811" number="8" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="2416" nation="BRA" region="PR" clubid="1404" swrid="93758" name="Apan/Maringá">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Isabel Henriques" birthdate="2007-09-05" gender="F" nation="BRA" license="414491" swrid="5755356" athleteid="1763" externalid="414491" level="MRGA">
              <RESULTS>
                <RESULT eventid="1077" points="140" swimtime="00:00:48.55" resultid="1764" heatid="4725" lane="4" entrytime="00:00:49.17" entrycourse="SCM" />
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="1765" heatid="4916" lane="4" />
                <RESULT eventid="1189" points="164" swimtime="00:01:31.78" resultid="1766" heatid="4936" lane="3" entrytime="00:01:30.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="188" swimtime="00:00:40.00" resultid="1767" heatid="5098" lane="3" entrytime="00:00:40.64" entrycourse="SCM" />
                <RESULT eventid="4417" points="136" swimtime="00:00:49.09" resultid="5676" heatid="4740" lane="4" />
                <RESULT eventid="5804" points="193" swimtime="00:00:39.65" resultid="10077" heatid="6063" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hammon" lastname="Henrique Costa" birthdate="2008-09-19" gender="M" nation="BRA" license="408703" swrid="5726000" athleteid="1756" externalid="408703" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="263" swimtime="00:00:33.93" resultid="1757" heatid="4785" lane="4" />
                <RESULT eventid="1105" points="242" swimtime="00:00:35.47" resultid="1758" heatid="4842" lane="2" />
                <RESULT eventid="1213" points="347" swimtime="00:01:18.66" resultid="1759" heatid="4955" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="332" swimtime="00:01:04.70" resultid="1760" heatid="5016" lane="4" entrytime="00:01:05.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="363" swimtime="00:00:28.26" resultid="1761" heatid="5224" lane="6" entrytime="00:00:28.73" entrycourse="SCM" />
                <RESULT eventid="1329" points="368" swimtime="00:00:34.79" resultid="1762" heatid="5157" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Garcia Cavalcante" birthdate="2011-11-21" gender="M" nation="BRA" license="378200" swrid="5603840" athleteid="1453" externalid="378200" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="211" swimtime="00:00:36.49" resultid="1454" heatid="4784" lane="2" />
                <RESULT eventid="1105" points="196" swimtime="00:00:38.02" resultid="1455" heatid="4843" lane="1" />
                <RESULT eventid="1213" points="302" swimtime="00:01:22.36" resultid="1456" heatid="4958" lane="2" entrytime="00:01:24.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="254" swimtime="00:03:09.61" resultid="1457" heatid="4995" lane="1" entrytime="00:03:06.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.71" />
                    <SPLIT distance="100" swimtime="00:01:30.49" />
                    <SPLIT distance="150" swimtime="00:02:20.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="264" swimtime="00:00:31.40" resultid="1458" heatid="5222" lane="3" entrytime="00:00:30.98" entrycourse="SCM" />
                <RESULT eventid="1329" points="252" swimtime="00:00:39.45" resultid="1459" heatid="5164" lane="1" entrytime="00:00:40.11" entrycourse="SCM" />
                <RESULT eventid="4429" points="187" swimtime="00:00:38.65" resultid="5762" heatid="4857" lane="6" />
                <RESULT eventid="5807" points="265" swimtime="00:00:38.80" resultid="10135" heatid="6041" lane="3" />
                <RESULT eventid="5810" points="267" swimtime="00:00:31.28" resultid="10251" heatid="6025" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Eduardo Ebiner" birthdate="2013-07-29" gender="M" nation="BRA" license="397371" swrid="5641763" athleteid="1689" externalid="397371" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="119" swimtime="00:00:44.20" resultid="1690" heatid="4786" lane="3" entrytime="00:00:46.76" entrycourse="SCM" />
                <RESULT eventid="1105" points="111" swimtime="00:00:45.94" resultid="1691" heatid="4847" lane="2" entrytime="00:00:48.18" entrycourse="SCM" />
                <RESULT eventid="1263" points="137" swimtime="00:03:52.97" resultid="1692" heatid="4994" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.00" />
                    <SPLIT distance="100" swimtime="00:01:52.07" />
                    <SPLIT distance="150" swimtime="00:02:53.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="147" swimtime="00:01:24.78" resultid="1693" heatid="5014" lane="5" entrytime="00:01:31.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="151" swimtime="00:00:37.85" resultid="1694" heatid="5217" lane="3" />
                <RESULT eventid="1329" points="121" swimtime="00:00:50.35" resultid="1695" heatid="5162" lane="3" entrytime="00:00:48.17" entrycourse="SCM" />
                <RESULT eventid="4423" points="121" swimtime="00:00:43.92" resultid="5697" heatid="4793" lane="4" />
                <RESULT eventid="4429" points="109" swimtime="00:00:46.18" resultid="5750" heatid="4853" lane="5" />
                <RESULT eventid="5807" points="123" swimtime="00:00:50.10" resultid="10125" heatid="6037" lane="4" />
                <RESULT eventid="5810" points="150" swimtime="00:00:37.94" resultid="10239" heatid="6021" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Donato De Morais" birthdate="2009-03-28" gender="F" nation="BRA" license="345588" swrid="5485198" athleteid="1516" externalid="345588" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="189" swimtime="00:00:42.45" resultid="1517" heatid="4673" lane="5" />
                <RESULT eventid="1077" points="248" swimtime="00:00:40.17" resultid="1518" heatid="4728" lane="3" entrytime="00:00:35.40" entrycourse="SCM" />
                <RESULT eventid="1119" status="DNS" swimtime="00:00:00.00" resultid="1519" heatid="4878" lane="3" entrytime="00:02:41.96" entrycourse="SCM" />
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="1520" heatid="4917" lane="3" entrytime="00:01:15.37" entrycourse="SCM" />
                <RESULT eventid="1314" points="238" swimtime="00:00:36.97" resultid="1521" heatid="5098" lane="6" />
                <RESULT eventid="1301" points="190" swimtime="00:00:49.30" resultid="1522" heatid="5048" lane="6" />
                <RESULT eventid="4411" points="191" swimtime="00:00:42.27" resultid="5629" heatid="4687" lane="2" />
                <RESULT eventid="4413" points="202" swimtime="00:00:41.51" resultid="5646" heatid="4694" lane="5" />
                <RESULT eventid="4417" points="262" swimtime="00:00:39.46" resultid="5671" heatid="4738" lane="1" />
                <RESULT eventid="4419" points="286" swimtime="00:00:38.32" resultid="5689" heatid="4745" lane="4" />
                <RESULT eventid="5801" points="183" swimtime="00:00:49.89" resultid="10034" heatid="6075" lane="2" />
                <RESULT eventid="5804" points="278" swimtime="00:00:35.13" resultid="10073" heatid="6061" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Pacheco" birthdate="2012-10-03" gender="M" nation="BRA" license="370663" swrid="5603883" athleteid="1551" externalid="370663" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="229" swimtime="00:00:35.50" resultid="1552" heatid="4789" lane="5" entrytime="00:00:34.37" entrycourse="SCM" />
                <RESULT eventid="1105" points="183" swimtime="00:00:38.90" resultid="1553" heatid="4849" lane="6" entrytime="00:00:40.43" entrycourse="SCM" />
                <RESULT eventid="1213" points="195" swimtime="00:01:35.28" resultid="1554" heatid="4958" lane="5" entrytime="00:01:33.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="259" swimtime="00:01:10.32" resultid="1555" heatid="5016" lane="6" entrytime="00:01:12.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="256" swimtime="00:00:31.72" resultid="1556" heatid="5222" lane="2" entrytime="00:00:31.96" entrycourse="SCM" />
                <RESULT eventid="1329" points="191" swimtime="00:00:43.31" resultid="1557" heatid="5163" lane="4" entrytime="00:00:43.64" entrycourse="SCM" />
                <RESULT eventid="4423" points="222" swimtime="00:00:35.87" resultid="5701" heatid="4795" lane="3" />
                <RESULT eventid="4429" points="159" swimtime="00:00:40.78" resultid="5756" heatid="4855" lane="6" />
                <RESULT eventid="5807" points="195" swimtime="00:00:43.02" resultid="10130" heatid="6039" lane="4" />
                <RESULT eventid="5810" points="253" swimtime="00:00:31.85" resultid="10243" heatid="6023" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Diogo" lastname="Sanchez" birthdate="2012-11-29" gender="M" nation="BRA" license="370658" swrid="5603906" athleteid="1425" externalid="370658" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="89" swimtime="00:00:48.59" resultid="1426" heatid="4786" lane="2" entrytime="00:00:53.33" entrycourse="SCM" />
                <RESULT eventid="1105" points="117" swimtime="00:00:45.14" resultid="1427" heatid="4848" lane="5" entrytime="00:00:44.69" entrycourse="SCM" />
                <RESULT eventid="1213" points="172" swimtime="00:01:39.40" resultid="1428" heatid="4957" lane="3" entrytime="00:01:42.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="162" swimtime="00:03:40.06" resultid="1429" heatid="4994" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.42" />
                    <SPLIT distance="100" swimtime="00:01:48.72" />
                    <SPLIT distance="150" swimtime="00:02:45.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="130" swimtime="00:00:39.78" resultid="1430" heatid="5220" lane="6" entrytime="00:00:36.70" entrycourse="SCM" />
                <RESULT eventid="1329" points="155" swimtime="00:00:46.38" resultid="1431" heatid="5163" lane="5" entrytime="00:00:44.88" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="De Desvars" birthdate="2016-04-08" gender="F" nation="BRA" license="414853" swrid="5757889" athleteid="1797" externalid="414853" level="MRGA">
              <RESULTS>
                <RESULT eventid="1117" points="56" swimtime="00:01:05.84" resultid="1798" heatid="4873" lane="4" entrytime="00:01:11.43" entrycourse="SCM" />
                <RESULT eventid="1141" points="28" swimtime="00:01:33.08" resultid="1799" heatid="4892" lane="4" entrytime="00:01:26.95" entrycourse="SCM" />
                <RESULT eventid="1177" points="42" swimtime="00:01:05.73" resultid="1800" heatid="4919" lane="4" entrytime="00:01:06.56" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Chaim" birthdate="2011-05-29" gender="F" nation="BRA" license="370662" swrid="5409721" athleteid="1488" externalid="370662" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="247" swimtime="00:00:38.84" resultid="1489" heatid="4675" lane="4" entrytime="00:00:42.81" entrycourse="SCM" />
                <RESULT eventid="1077" points="246" swimtime="00:00:40.28" resultid="1490" heatid="4727" lane="6" entrytime="00:00:41.38" entrycourse="SCM" />
                <RESULT eventid="1143" points="324" swimtime="00:02:40.54" resultid="1491" heatid="4897" lane="1" entrytime="00:02:41.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                    <SPLIT distance="100" swimtime="00:01:16.91" />
                    <SPLIT distance="150" swimtime="00:01:59.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="336" swimtime="00:01:12.28" resultid="1492" heatid="4938" lane="4" entrytime="00:01:13.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="241" swimtime="00:00:36.82" resultid="1493" heatid="5101" lane="3" entrytime="00:00:33.57" entrycourse="SCM" />
                <RESULT eventid="1301" points="213" swimtime="00:00:47.46" resultid="1494" heatid="5047" lane="4" />
                <RESULT eventid="4411" points="247" swimtime="00:00:38.85" resultid="5620" heatid="4683" lane="2" />
                <RESULT eventid="4413" points="228" swimtime="00:00:39.88" resultid="5640" heatid="4692" lane="5" />
                <RESULT eventid="4417" points="250" swimtime="00:00:40.03" resultid="5662" heatid="4734" lane="1" />
                <RESULT eventid="4419" points="277" swimtime="00:00:38.73" resultid="5684" heatid="4743" lane="5" />
                <RESULT eventid="5801" points="203" swimtime="00:00:48.27" resultid="10024" heatid="6071" lane="2" />
                <RESULT eventid="5804" points="342" swimtime="00:00:32.76" resultid="10066" heatid="6057" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolas" lastname="Baldo De França" birthdate="2014-04-21" gender="M" nation="BRA" license="393773" swrid="5507467" athleteid="1661" externalid="393773" level="MRGA">
              <RESULTS>
                <RESULT eventid="1089" points="99" swimtime="00:00:46.86" resultid="1662" heatid="4759" lane="2" entrytime="00:00:48.49" entrycourse="SCM" />
                <RESULT eventid="1102" points="57" swimtime="00:00:57.26" resultid="1663" heatid="4818" lane="3" />
                <RESULT eventid="1213" points="83" swimtime="00:02:06.56" resultid="1664" heatid="4955" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="84" swimtime="00:01:42.11" resultid="1665" heatid="5013" lane="1" entrytime="00:01:39.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="107" swimtime="00:00:42.43" resultid="1666" heatid="5192" lane="3" entrytime="00:00:45.96" entrycourse="SCM" />
                <RESULT eventid="1326" points="86" swimtime="00:00:56.48" resultid="1667" heatid="5133" lane="1" entrytime="00:00:58.02" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Vaneti Mazuti" birthdate="2014-11-29" gender="M" nation="BRA" license="414850" swrid="5757897" athleteid="1779" externalid="414850" level="MRGA">
              <RESULTS>
                <RESULT eventid="1089" status="DNS" swimtime="00:00:00.00" resultid="1780" heatid="4758" lane="3" entrytime="00:00:55.94" entrycourse="SCM" />
                <RESULT eventid="1102" status="DNS" swimtime="00:00:00.00" resultid="1781" heatid="4818" lane="5" />
                <RESULT eventid="1213" status="DNS" swimtime="00:00:00.00" resultid="1782" heatid="4957" lane="5" />
                <RESULT eventid="1249" status="DNS" swimtime="00:00:00.00" resultid="1783" heatid="4987" lane="4" />
                <RESULT eventid="1285" status="DNS" swimtime="00:00:00.00" resultid="1784" heatid="5192" lane="4" entrytime="00:00:46.13" entrycourse="SCM" />
                <RESULT eventid="1326" status="DNS" swimtime="00:00:00.00" resultid="1785" heatid="5134" lane="2" entrytime="00:00:51.55" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio" lastname="Rafael Padial" birthdate="2014-03-07" gender="M" nation="BRA" license="397331" swrid="5641774" athleteid="1682" externalid="397331" level="MRGA">
              <RESULTS>
                <RESULT eventid="1089" points="116" swimtime="00:00:44.56" resultid="1683" heatid="4759" lane="4" entrytime="00:00:44.98" entrycourse="SCM" />
                <RESULT eventid="1102" points="121" swimtime="00:00:44.59" resultid="1684" heatid="4820" lane="3" entrytime="00:00:42.10" entrycourse="SCM" />
                <RESULT eventid="1249" points="129" swimtime="00:01:35.42" resultid="1685" heatid="4988" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="159" swimtime="00:01:22.75" resultid="1686" heatid="5015" lane="1" entrytime="00:01:20.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="179" swimtime="00:00:35.74" resultid="1687" heatid="5194" lane="4" entrytime="00:00:35.06" entrycourse="SCM" />
                <RESULT eventid="1326" points="130" swimtime="00:00:49.14" resultid="1688" heatid="5134" lane="5" entrytime="00:00:51.83" entrycourse="SCM" />
                <RESULT eventid="4421" points="111" swimtime="00:00:45.18" resultid="9027" heatid="9006" lane="6" />
                <RESULT eventid="4427" points="124" swimtime="00:00:44.27" resultid="9032" heatid="9008" lane="5" />
                <RESULT eventid="4445" points="123" swimtime="00:00:50.15" resultid="10118" heatid="6035" lane="3" />
                <RESULT eventid="4451" points="180" swimtime="00:00:35.64" resultid="10230" heatid="6019" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Rampasi" birthdate="2013-10-16" gender="F" nation="BRA" license="382209" swrid="5603866" athleteid="1605" externalid="382209" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="114" swimtime="00:00:50.24" resultid="1606" heatid="4675" lane="6" entrytime="00:00:48.10" entrycourse="SCM" />
                <RESULT eventid="1077" points="112" swimtime="00:00:52.30" resultid="1607" heatid="4725" lane="5" entrytime="00:00:53.42" entrycourse="SCM" />
                <RESULT eventid="1143" points="219" swimtime="00:03:02.88" resultid="1608" heatid="4896" lane="4" entrytime="00:03:09.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.35" />
                    <SPLIT distance="100" swimtime="00:01:33.18" />
                    <SPLIT distance="150" swimtime="00:02:19.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="194" swimtime="00:01:26.72" resultid="1609" heatid="4937" lane="6" entrytime="00:01:30.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="191" swimtime="00:00:39.77" resultid="1610" heatid="5099" lane="6" entrytime="00:00:39.88" entrycourse="SCM" />
                <RESULT eventid="1301" points="135" swimtime="00:00:55.26" resultid="1611" heatid="5049" lane="1" entrytime="00:00:55.36" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Muniz" birthdate="2012-09-03" gender="M" nation="BRA" license="392106" swrid="5603877" athleteid="1633" externalid="392106" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="128" swimtime="00:00:43.13" resultid="1634" heatid="4787" lane="6" entrytime="00:00:46.42" entrycourse="SCM" />
                <RESULT eventid="1105" points="127" swimtime="00:00:43.91" resultid="1635" heatid="4847" lane="4" entrytime="00:00:47.51" entrycourse="SCM" />
                <RESULT eventid="1227" points="186" swimtime="00:02:53.94" resultid="1636" heatid="4968" lane="3" entrytime="00:03:06.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.72" />
                    <SPLIT distance="100" swimtime="00:01:24.61" />
                    <SPLIT distance="150" swimtime="00:02:10.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="196" swimtime="00:01:17.15" resultid="1637" heatid="5015" lane="6" entrytime="00:01:21.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="207" swimtime="00:00:34.03" resultid="1638" heatid="5220" lane="4" entrytime="00:00:35.40" entrycourse="SCM" />
                <RESULT eventid="1329" points="119" swimtime="00:00:50.72" resultid="1639" heatid="5160" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sara" lastname="Padovin Chiste" birthdate="2015-02-04" gender="F" nation="BRA" license="414849" swrid="5755358" athleteid="1772" externalid="414849" level="MRGA">
              <RESULTS>
                <RESULT eventid="1061" status="DNS" swimtime="00:00:00.00" resultid="1773" heatid="4653" lane="3" entrytime="00:01:05.81" entrycourse="SCM" />
                <RESULT eventid="1074" status="DNS" swimtime="00:00:00.00" resultid="1774" heatid="4703" lane="4" />
                <RESULT eventid="1129" points="123" swimtime="00:02:05.22" resultid="1775" heatid="4889" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="99" swimtime="00:01:48.31" resultid="1776" heatid="4936" lane="6" entrytime="00:01:51.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="107" swimtime="00:00:59.71" resultid="1777" heatid="5027" lane="4" entrytime="00:01:00.75" entrycourse="SCM" />
                <RESULT eventid="1311" points="90" swimtime="00:00:50.98" resultid="1778" heatid="5077" lane="4" entrytime="00:00:53.44" entrycourse="SCM" />
                <RESULT eventid="4433" points="109" swimtime="00:00:59.34" resultid="10001" heatid="5030" lane="1" />
                <RESULT eventid="4439" points="102" swimtime="00:00:48.98" resultid="10039" heatid="6049" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felype" lastname="Gongora Zago" birthdate="2011-09-14" gender="M" nation="BRA" license="392099" swrid="5603848" athleteid="1460" externalid="392099" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="254" swimtime="00:00:34.30" resultid="1461" heatid="4788" lane="4" entrytime="00:00:35.97" entrycourse="SCM" />
                <RESULT eventid="1105" points="181" swimtime="00:00:39.05" resultid="1462" heatid="4842" lane="3" />
                <RESULT eventid="1203" points="199" swimtime="00:03:00.87" resultid="1463" heatid="4944" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.87" />
                    <SPLIT distance="100" swimtime="00:01:28.21" />
                    <SPLIT distance="150" swimtime="00:02:16.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="242" swimtime="00:01:11.94" resultid="1464" heatid="5015" lane="4" entrytime="00:01:14.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="247" swimtime="00:00:32.13" resultid="1465" heatid="5221" lane="4" entrytime="00:00:33.10" entrycourse="SCM" />
                <RESULT eventid="1329" points="141" swimtime="00:00:47.92" resultid="1466" heatid="5161" lane="1" />
                <RESULT eventid="4423" points="214" swimtime="00:00:36.35" resultid="5710" heatid="4797" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Campos" birthdate="2013-02-17" gender="M" nation="BRA" license="377262" swrid="5641756" athleteid="1579" externalid="377262" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="106" swimtime="00:00:45.95" resultid="1580" heatid="4787" lane="5" entrytime="00:00:44.99" entrycourse="SCM" />
                <RESULT eventid="1105" points="150" swimtime="00:00:41.53" resultid="1581" heatid="4849" lane="5" entrytime="00:00:39.51" entrycourse="SCM" />
                <RESULT eventid="1227" points="188" swimtime="00:02:53.22" resultid="1582" heatid="5254" lane="5" entrytime="00:02:59.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.95" />
                    <SPLIT distance="100" swimtime="00:01:26.12" />
                    <SPLIT distance="150" swimtime="00:02:10.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="151" swimtime="00:01:30.66" resultid="1583" heatid="4988" lane="2" entrytime="00:01:27.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="185" swimtime="00:00:35.34" resultid="1584" heatid="5220" lane="1" entrytime="00:00:36.40" entrycourse="SCM" />
                <RESULT eventid="1329" points="113" swimtime="00:00:51.51" resultid="1585" heatid="5159" lane="1" />
                <RESULT eventid="4423" points="113" swimtime="00:00:44.89" resultid="5698" heatid="4793" lane="5" />
                <RESULT eventid="4429" points="155" swimtime="00:00:41.14" resultid="5746" heatid="4853" lane="1" />
                <RESULT eventid="4431" points="161" swimtime="00:00:40.56" resultid="5777" heatid="4864" lane="4" />
                <RESULT eventid="5807" points="114" swimtime="00:00:51.31" resultid="10126" heatid="6037" lane="5" />
                <RESULT eventid="5810" points="187" swimtime="00:00:35.25" resultid="10238" heatid="6021" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnes" lastname="Sophie Amadei" birthdate="2014-01-10" gender="F" nation="BRA" license="403388" swrid="5676293" athleteid="1715" externalid="403388" level="MRGA">
              <RESULTS>
                <RESULT eventid="1061" points="108" swimtime="00:00:51.13" resultid="1716" heatid="4654" lane="5" entrytime="00:00:52.80" entrycourse="SCM" />
                <RESULT eventid="1074" points="87" swimtime="00:00:56.96" resultid="1717" heatid="4704" lane="2" entrytime="00:01:04.08" entrycourse="SCM" />
                <RESULT eventid="1129" points="113" swimtime="00:02:08.63" resultid="1718" heatid="4888" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" status="DNS" swimtime="00:00:00.00" resultid="1719" heatid="4902" lane="3" />
                <RESULT eventid="1298" points="113" swimtime="00:00:58.54" resultid="1720" heatid="5027" lane="3" entrytime="00:00:58.73" entrycourse="SCM" />
                <RESULT eventid="1311" points="155" swimtime="00:00:42.64" resultid="1721" heatid="5078" lane="2" entrytime="00:00:45.81" entrycourse="SCM" />
                <RESULT eventid="4439" points="163" swimtime="00:00:41.94" resultid="10049" heatid="6051" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raphael" lastname="Piai Pellegrini" birthdate="2012-03-24" gender="M" nation="BRA" license="377261" swrid="5603894" athleteid="1572" externalid="377261" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="294" swimtime="00:00:32.68" resultid="1573" heatid="4789" lane="4" entrytime="00:00:32.95" entrycourse="SCM" />
                <RESULT eventid="1105" points="197" swimtime="00:00:37.96" resultid="1574" heatid="4849" lane="4" entrytime="00:00:35.58" entrycourse="SCM" />
                <RESULT eventid="1237" points="261" swimtime="00:01:14.69" resultid="1575" heatid="4976" lane="2" entrytime="00:01:15.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="331" swimtime="00:01:04.81" resultid="1576" heatid="5017" lane="6" entrytime="00:01:04.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="248" swimtime="00:00:32.07" resultid="1577" heatid="5223" lane="3" entrytime="00:00:29.00" entrycourse="SCM" />
                <RESULT eventid="1329" points="215" swimtime="00:00:41.62" resultid="1578" heatid="5161" lane="2" />
                <RESULT eventid="4423" points="299" swimtime="00:00:32.52" resultid="5699" heatid="4795" lane="1" />
                <RESULT eventid="4425" points="309" swimtime="00:00:32.16" resultid="5731" heatid="4805" lane="4" />
                <RESULT eventid="4429" points="181" swimtime="00:00:39.02" resultid="5754" heatid="4855" lane="4" />
                <RESULT eventid="5807" points="225" swimtime="00:00:41.01" resultid="10128" heatid="6039" lane="2" />
                <RESULT eventid="5810" points="336" swimtime="00:00:28.98" resultid="10244" heatid="6023" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="De Correa" birthdate="2014-12-03" gender="M" nation="BRA" license="403387" swrid="5676286" athleteid="1708" externalid="403387" level="MRGA">
              <RESULTS>
                <RESULT eventid="1089" points="132" swimtime="00:00:42.64" resultid="1709" heatid="4757" lane="5" />
                <RESULT eventid="1102" points="98" swimtime="00:00:47.88" resultid="1710" heatid="4820" lane="5" entrytime="00:00:46.16" entrycourse="SCM" />
                <RESULT eventid="1249" points="99" swimtime="00:01:44.20" resultid="1711" heatid="4988" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="128" swimtime="00:01:28.89" resultid="1712" heatid="5014" lane="1" entrytime="00:01:32.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="142" swimtime="00:00:38.57" resultid="1713" heatid="5194" lane="1" entrytime="00:00:39.33" entrycourse="SCM" />
                <RESULT eventid="1326" points="91" swimtime="00:00:55.38" resultid="1714" heatid="5133" lane="2" entrytime="00:00:56.43" entrycourse="SCM" />
                <RESULT eventid="4421" points="127" swimtime="00:00:43.20" resultid="9026" heatid="9006" lane="5" />
                <RESULT eventid="4445" points="91" swimtime="00:00:55.45" resultid="10121" heatid="6035" lane="6" />
                <RESULT eventid="4451" points="143" swimtime="00:00:38.51" resultid="10231" heatid="6019" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Otavio Luz" birthdate="2013-07-27" gender="M" nation="BRA" license="392111" swrid="5603882" athleteid="1654" externalid="392111" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="185" swimtime="00:00:38.11" resultid="1655" heatid="4787" lane="4" entrytime="00:00:39.22" entrycourse="SCM" />
                <RESULT eventid="1105" points="144" swimtime="00:00:42.15" resultid="1656" heatid="4848" lane="6" entrytime="00:00:45.05" entrycourse="SCM" />
                <RESULT eventid="1203" points="151" swimtime="00:03:18.00" resultid="1657" heatid="4945" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.52" />
                    <SPLIT distance="100" swimtime="00:01:38.55" />
                    <SPLIT distance="150" swimtime="00:02:30.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1237" points="156" swimtime="00:01:28.70" resultid="1658" heatid="4976" lane="5" entrytime="00:01:28.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="200" swimtime="00:00:34.47" resultid="1659" heatid="5220" lane="2" entrytime="00:00:35.59" entrycourse="SCM" />
                <RESULT eventid="1329" points="140" swimtime="00:00:48.05" resultid="1660" heatid="5162" lane="2" entrytime="00:00:49.95" entrycourse="SCM" />
                <RESULT eventid="4423" points="176" swimtime="00:00:38.77" resultid="5694" heatid="4793" lane="1" />
                <RESULT eventid="4425" points="184" swimtime="00:00:38.22" resultid="5728" heatid="4804" lane="4" />
                <RESULT eventid="4429" points="149" swimtime="00:00:41.70" resultid="5747" heatid="4853" lane="2" />
                <RESULT eventid="4431" points="160" swimtime="00:00:40.69" resultid="5779" heatid="4864" lane="6" />
                <RESULT eventid="5807" points="136" swimtime="00:00:48.47" resultid="10123" heatid="6037" lane="2" />
                <RESULT eventid="5810" points="202" swimtime="00:00:34.34" resultid="10235" heatid="6021" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Pacheco" birthdate="2006-12-20" gender="M" nation="BRA" license="336850" swrid="5603854" athleteid="1502" externalid="336850" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="449" swimtime="00:00:28.40" resultid="1503" heatid="4791" lane="6" entrytime="00:00:28.63" entrycourse="SCM" />
                <RESULT eventid="1105" points="356" swimtime="00:00:31.18" resultid="1504" heatid="4845" lane="2" />
                <RESULT eventid="1237" points="398" swimtime="00:01:04.94" resultid="1505" heatid="4977" lane="5" entrytime="00:01:02.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="437" swimtime="00:00:59.05" resultid="1506" heatid="5018" lane="5" entrytime="00:00:56.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="1507" heatid="5218" lane="3" />
                <RESULT eventid="1329" status="DNS" swimtime="00:00:00.00" resultid="1508" heatid="5161" lane="4" />
                <RESULT eventid="4423" points="426" swimtime="00:00:28.89" resultid="5724" heatid="4803" lane="4" />
                <RESULT eventid="4429" points="345" swimtime="00:00:31.51" resultid="5775" heatid="4863" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Campelo" birthdate="2011-09-12" gender="M" nation="BRA" license="366963" swrid="5588742" athleteid="1405" externalid="366963" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="379" swimtime="00:00:30.05" resultid="1406" heatid="4790" lane="1" entrytime="00:00:30.43" entrycourse="SCM" />
                <RESULT eventid="1105" points="271" swimtime="00:00:34.15" resultid="1407" heatid="4851" lane="6" entrytime="00:00:30.81" entrycourse="SCM" />
                <RESULT eventid="1227" points="422" swimtime="00:02:12.41" resultid="1408" heatid="5254" lane="4" entrytime="00:02:21.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.02" />
                    <SPLIT distance="100" swimtime="00:01:06.22" />
                    <SPLIT distance="150" swimtime="00:01:40.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="449" swimtime="00:00:58.52" resultid="1409" heatid="5018" lane="6" entrytime="00:00:58.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="363" swimtime="00:00:28.26" resultid="1410" heatid="5225" lane="3" entrytime="00:00:26.31" entrycourse="SCM" />
                <RESULT eventid="1329" points="292" swimtime="00:00:37.59" resultid="1411" heatid="5158" lane="4" />
                <RESULT eventid="4423" points="313" swimtime="00:00:32.01" resultid="5705" heatid="4797" lane="1" />
                <RESULT eventid="4425" points="423" swimtime="00:00:28.96" resultid="5736" heatid="4806" lane="6" />
                <RESULT eventid="4429" points="285" swimtime="00:00:33.56" resultid="5758" heatid="4857" lane="2" />
                <RESULT eventid="4431" points="404" swimtime="00:00:29.89" resultid="5784" heatid="4866" lane="5" />
                <RESULT eventid="5807" points="320" swimtime="00:00:36.46" resultid="10133" heatid="6041" lane="1" />
                <RESULT eventid="5810" points="473" swimtime="00:00:25.86" resultid="10246" heatid="6025" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wellington" lastname="De Lima" birthdate="2008-03-01" gender="M" nation="BRA" license="370024" swrid="5470912" athleteid="1432" externalid="370024" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="446" swimtime="00:00:28.46" resultid="1433" heatid="4785" lane="5" />
                <RESULT eventid="1105" points="387" swimtime="00:00:30.32" resultid="1434" heatid="4851" lane="1" entrytime="00:00:30.25" entrycourse="SCM" />
                <RESULT eventid="1227" points="493" swimtime="00:02:05.72" resultid="1435" heatid="4968" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.46" />
                    <SPLIT distance="100" swimtime="00:01:00.26" />
                    <SPLIT distance="150" swimtime="00:01:33.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="485" swimtime="00:00:57.04" resultid="1436" heatid="5018" lane="2" entrytime="00:00:56.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="452" swimtime="00:00:26.26" resultid="1437" heatid="5226" lane="6" entrytime="00:00:25.87" entrycourse="SCM" />
                <RESULT eventid="1329" points="395" swimtime="00:00:33.99" resultid="1438" heatid="5156" lane="3" />
                <RESULT eventid="4423" points="439" swimtime="00:00:28.60" resultid="5726" heatid="4803" lane="5" />
                <RESULT eventid="4425" points="425" swimtime="00:00:28.92" resultid="5745" heatid="4809" lane="6" />
                <RESULT eventid="4429" points="414" swimtime="00:00:29.66" resultid="5774" heatid="4863" lane="4" />
                <RESULT eventid="5810" points="451" swimtime="00:00:26.27" resultid="10266" heatid="6031" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Antonio Mendes" birthdate="2008-12-04" gender="M" nation="BRA" license="366962" swrid="5196287" athleteid="1530" externalid="366962" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="438" swimtime="00:00:28.63" resultid="1531" heatid="4786" lane="1" />
                <RESULT eventid="1105" points="418" swimtime="00:00:29.56" resultid="1532" heatid="4851" lane="5" entrytime="00:00:30.20" entrycourse="SCM" />
                <RESULT eventid="1203" points="431" swimtime="00:02:19.74" resultid="1533" heatid="4945" lane="3" entrytime="00:02:25.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                    <SPLIT distance="100" swimtime="00:01:07.04" />
                    <SPLIT distance="150" swimtime="00:01:43.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="527" swimtime="00:01:08.40" resultid="1534" heatid="4959" lane="4" entrytime="00:01:08.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="419" swimtime="00:00:26.94" resultid="1535" heatid="5225" lane="2" entrytime="00:00:26.95" entrycourse="SCM" />
                <RESULT eventid="1329" points="478" swimtime="00:00:31.89" resultid="1536" heatid="5165" lane="4" entrytime="00:00:31.32" entrycourse="SCM" />
                <RESULT eventid="4429" points="421" swimtime="00:00:29.50" resultid="5773" heatid="4863" lane="3" />
                <RESULT eventid="4431" points="402" swimtime="00:00:29.95" resultid="5794" heatid="4869" lane="6" />
                <RESULT eventid="5807" points="506" swimtime="00:00:31.31" resultid="10151" heatid="6047" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Marques" birthdate="2015-10-15" gender="F" nation="BRA" license="399738" swrid="5651346" athleteid="1703" externalid="399738" level="MRGA">
              <RESULTS>
                <RESULT eventid="1061" points="20" swimtime="00:01:29.26" resultid="1704" heatid="4652" lane="5" />
                <RESULT eventid="1074" points="49" swimtime="00:01:08.94" resultid="1705" heatid="4704" lane="5" entrytime="00:01:08.91" entrycourse="SCM" />
                <RESULT eventid="1298" points="29" swimtime="00:01:31.86" resultid="1706" heatid="5026" lane="3" entrytime="00:01:35.58" entrycourse="SCM" />
                <RESULT eventid="1311" points="39" swimtime="00:01:07.55" resultid="1707" heatid="5077" lane="5" entrytime="00:01:12.64" entrycourse="SCM" />
                <RESULT eventid="4415" points="44" swimtime="00:01:11.37" resultid="9011" heatid="9003" lane="5" />
                <RESULT eventid="4409" points="14" swimtime="00:01:40.47" resultid="9017" heatid="9001" lane="6" />
                <RESULT eventid="4433" points="36" swimtime="00:01:25.33" resultid="10004" heatid="5030" lane="4" />
                <RESULT eventid="4439" points="45" swimtime="00:01:04.05" resultid="10043" heatid="6049" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Peroni Passafaro" birthdate="2013-09-17" gender="F" nation="BRA" license="370659" swrid="5603893" athleteid="1544" externalid="370659" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" status="DNS" swimtime="00:00:00.00" resultid="1545" heatid="4676" lane="1" entrytime="00:00:40.41" entrycourse="SCM" />
                <RESULT eventid="1077" status="DNS" swimtime="00:00:00.00" resultid="1546" heatid="4726" lane="5" entrytime="00:00:45.15" entrycourse="SCM" />
                <RESULT eventid="1119" status="DNS" swimtime="00:00:00.00" resultid="1547" heatid="4878" lane="2" />
                <RESULT eventid="1189" status="DNS" swimtime="00:00:00.00" resultid="1548" heatid="4939" lane="6" entrytime="00:01:20.44" entrycourse="SCM" />
                <RESULT eventid="1314" status="DNS" swimtime="00:00:00.00" resultid="1549" heatid="5100" lane="2" entrytime="00:00:35.21" entrycourse="SCM" />
                <RESULT eventid="1301" status="DNS" swimtime="00:00:00.00" resultid="1550" heatid="5047" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Coleto Arcanjo" birthdate="2015-08-17" gender="F" nation="BRA" license="407176" swrid="5631404" athleteid="1734" externalid="407176" level="MRGA">
              <RESULTS>
                <RESULT eventid="1061" points="29" swimtime="00:01:18.82" resultid="1735" heatid="4653" lane="4" entrytime="00:01:17.90" entrycourse="SCM" />
                <RESULT eventid="1074" points="46" swimtime="00:01:10.29" resultid="1736" heatid="4704" lane="1" entrytime="00:01:13.77" entrycourse="SCM" />
                <RESULT eventid="1298" points="46" swimtime="00:01:19.02" resultid="1737" heatid="5027" lane="6" entrytime="00:01:18.10" entrycourse="SCM" />
                <RESULT eventid="1311" points="43" swimtime="00:01:05.45" resultid="1738" heatid="5077" lane="2" entrytime="00:01:07.66" entrycourse="SCM" />
                <RESULT eventid="4415" points="52" swimtime="00:01:07.52" resultid="9010" heatid="9003" lane="6" />
                <RESULT eventid="4409" points="25" swimtime="00:01:23.27" resultid="9016" heatid="9001" lane="5" />
                <RESULT eventid="4433" points="32" swimtime="00:01:28.55" resultid="10003" heatid="5030" lane="3" />
                <RESULT eventid="4439" points="45" swimtime="00:01:04.15" resultid="10042" heatid="6049" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Forti Francisco" birthdate="2015-07-08" gender="M" nation="BRA" license="392104" swrid="5534395" athleteid="1626" externalid="392104" level="MRGA">
              <RESULTS>
                <RESULT eventid="1089" points="70" swimtime="00:00:52.76" resultid="1627" heatid="4758" lane="4" entrytime="00:00:57.51" entrycourse="SCM" />
                <RESULT eventid="1102" points="72" swimtime="00:00:53.03" resultid="1628" heatid="4818" lane="4" />
                <RESULT eventid="1213" points="93" swimtime="00:02:01.73" resultid="1629" heatid="4956" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="93" swimtime="00:01:38.88" resultid="1630" heatid="5014" lane="6" entrytime="00:01:33.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" status="DNS" swimtime="00:00:00.00" resultid="1631" heatid="5194" lane="6" entrytime="00:00:41.32" entrycourse="SCM" />
                <RESULT eventid="1326" status="DNS" swimtime="00:00:00.00" resultid="1632" heatid="5133" lane="4" entrytime="00:00:56.39" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Quental De Meireles" birthdate="2008-11-20" gender="M" nation="BRA" license="392103" swrid="5603898" athleteid="1474" externalid="392103" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="378" swimtime="00:00:30.07" resultid="1475" heatid="4790" lane="2" entrytime="00:00:30.24" entrycourse="SCM" />
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="1476" heatid="4845" lane="5" />
                <RESULT eventid="1237" status="DNS" swimtime="00:00:00.00" resultid="1477" heatid="4977" lane="6" entrytime="00:01:07.49" entrycourse="SCM" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="1478" heatid="5017" lane="1" entrytime="00:01:04.27" entrycourse="SCM" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="1479" heatid="5224" lane="4" entrytime="00:00:28.38" entrycourse="SCM" />
                <RESULT eventid="1329" status="DNS" swimtime="00:00:00.00" resultid="1480" heatid="5159" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Bessa" birthdate="2003-06-19" gender="M" nation="BRA" license="317841" swrid="5312237" athleteid="1412" externalid="317841" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="425" swimtime="00:00:28.91" resultid="1413" heatid="4786" lane="6" />
                <RESULT eventid="1105" points="332" swimtime="00:00:31.91" resultid="1414" heatid="4844" lane="4" />
                <RESULT eventid="1213" points="620" swimtime="00:01:04.82" resultid="1415" heatid="4959" lane="3" entrytime="00:01:04.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="454" swimtime="00:00:26.23" resultid="1416" heatid="5226" lane="1" entrytime="00:00:25.28" entrycourse="SCM" />
                <RESULT eventid="1329" points="534" swimtime="00:00:30.74" resultid="1417" heatid="5165" lane="3" entrytime="00:00:29.77" entrycourse="SCM" />
                <RESULT eventid="4429" points="355" swimtime="00:00:31.22" resultid="5776" heatid="4863" lane="6" />
                <RESULT eventid="5807" points="583" swimtime="00:00:29.86" resultid="10149" heatid="6047" lane="2" />
                <RESULT eventid="5810" points="402" swimtime="00:00:27.31" resultid="10265" heatid="6031" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Ghelere" birthdate="2011-04-03" gender="F" nation="BRA" license="368146" swrid="5603843" athleteid="1495" externalid="368146" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="300" swimtime="00:00:36.39" resultid="1496" heatid="4672" lane="4" />
                <RESULT eventid="1077" points="221" swimtime="00:00:41.75" resultid="1497" heatid="4724" lane="5" />
                <RESULT eventid="1153" points="195" swimtime="00:01:33.17" resultid="1498" heatid="4903" lane="1" entrytime="00:01:28.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="282" swimtime="00:01:16.62" resultid="1499" heatid="4938" lane="3" entrytime="00:01:10.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="271" swimtime="00:00:35.43" resultid="1500" heatid="5102" lane="4" entrytime="00:00:32.30" entrycourse="SCM" />
                <RESULT eventid="1301" points="171" swimtime="00:00:51.02" resultid="1501" heatid="5049" lane="6" />
                <RESULT eventid="4411" points="259" swimtime="00:00:38.21" resultid="5619" heatid="4683" lane="1" />
                <RESULT eventid="4413" points="305" swimtime="00:00:36.18" resultid="5639" heatid="4692" lane="4" />
                <RESULT eventid="4417" points="252" swimtime="00:00:39.96" resultid="5664" heatid="4734" lane="3" />
                <RESULT eventid="4419" points="276" swimtime="00:00:38.78" resultid="5683" heatid="4743" lane="4" />
                <RESULT comment="SW 7.1 - Mais de uma pernada de borboleta antes da primeira pernada de peito após o início ou a virada.  (Horário: 9:54), Após a volta dos 25m." eventid="5801" status="DSQ" swimtime="00:00:49.88" resultid="10026" heatid="6071" lane="4" />
                <RESULT eventid="5804" points="279" swimtime="00:00:35.05" resultid="10064" heatid="6057" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lara" lastname="Constantino" birthdate="2012-06-02" gender="F" nation="BRA" license="382208" swrid="5420069" athleteid="1598" externalid="382208" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="232" swimtime="00:00:39.66" resultid="1599" heatid="4676" lane="5" entrytime="00:00:40.31" entrycourse="SCM" />
                <RESULT eventid="1077" points="184" swimtime="00:00:44.32" resultid="1600" heatid="4727" lane="1" entrytime="00:00:41.10" entrycourse="SCM" />
                <RESULT eventid="1129" points="315" swimtime="00:01:31.56" resultid="1601" heatid="4890" lane="1" entrytime="00:01:37.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="279" swimtime="00:03:25.70" resultid="1602" heatid="4923" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.94" />
                    <SPLIT distance="100" swimtime="00:01:40.37" />
                    <SPLIT distance="150" swimtime="00:02:34.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="244" swimtime="00:00:36.65" resultid="1603" heatid="5102" lane="1" entrytime="00:00:33.31" entrycourse="SCM" />
                <RESULT eventid="1301" points="293" swimtime="00:00:42.71" resultid="1604" heatid="5051" lane="1" entrytime="00:00:41.26" entrycourse="SCM" />
                <RESULT eventid="4411" points="196" swimtime="00:00:41.91" resultid="5617" heatid="4681" lane="5" />
                <RESULT eventid="4417" points="194" swimtime="00:00:43.60" resultid="5661" heatid="4732" lane="6" />
                <RESULT eventid="5801" points="301" swimtime="00:00:42.29" resultid="10020" heatid="6069" lane="4" />
                <RESULT eventid="5804" points="297" swimtime="00:00:34.33" resultid="10060" heatid="6055" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Garcia Cavalcante" birthdate="2008-08-11" gender="M" nation="BRA" license="369676" swrid="5603841" athleteid="1446" externalid="369676" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="291" swimtime="00:00:32.81" resultid="1447" heatid="4784" lane="5" />
                <RESULT eventid="1105" points="240" swimtime="00:00:35.54" resultid="1448" heatid="4846" lane="5" />
                <RESULT eventid="1263" points="417" swimtime="00:02:40.78" resultid="1449" heatid="4995" lane="2" entrytime="00:02:41.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.46" />
                    <SPLIT distance="100" swimtime="00:01:17.52" />
                    <SPLIT distance="150" swimtime="00:01:58.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="368" swimtime="00:01:02.56" resultid="1450" heatid="5017" lane="2" entrytime="00:01:00.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="328" swimtime="00:00:29.22" resultid="1451" heatid="5224" lane="2" entrytime="00:00:28.39" entrycourse="SCM" />
                <RESULT eventid="1329" points="383" swimtime="00:00:34.33" resultid="1452" heatid="5160" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laion" lastname="Miguel Simoes" birthdate="2016-04-02" gender="M" nation="BRA" license="407179" swrid="5718695" athleteid="1739" externalid="407179" level="MRGA">
              <RESULTS>
                <RESULT eventid="1201" points="71" swimtime="00:00:53.32" resultid="1740" heatid="4941" lane="2" entrytime="00:01:02.90" entrycourse="SCM" />
                <RESULT eventid="1225" points="62" swimtime="00:01:02.99" resultid="1741" heatid="4961" lane="4" entrytime="00:01:05.42" entrycourse="SCM" />
                <RESULT eventid="1261" points="100" swimtime="00:00:43.43" resultid="1742" heatid="4991" lane="2" entrytime="00:00:50.58" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Tomazeli" birthdate="2013-02-05" gender="M" nation="BRA" license="392109" swrid="5614097" athleteid="1647" externalid="392109" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="148" swimtime="00:00:41.08" resultid="1648" heatid="4787" lane="2" entrytime="00:00:44.06" entrycourse="SCM" />
                <RESULT eventid="1105" points="127" swimtime="00:00:43.96" resultid="1649" heatid="4848" lane="2" entrytime="00:00:44.00" entrycourse="SCM" />
                <RESULT eventid="1227" points="180" swimtime="00:02:55.69" resultid="1650" heatid="5254" lane="6" entrytime="00:03:03.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.77" />
                    <SPLIT distance="100" swimtime="00:01:27.70" />
                    <SPLIT distance="150" swimtime="00:02:13.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1237" points="101" swimtime="00:01:42.56" resultid="1651" heatid="4977" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="191" swimtime="00:00:34.99" resultid="1652" heatid="5219" lane="3" entrytime="00:00:36.82" entrycourse="SCM" />
                <RESULT eventid="1329" points="123" swimtime="00:00:50.15" resultid="1653" heatid="5162" lane="1" entrytime="00:00:51.89" entrycourse="SCM" />
                <RESULT eventid="4423" points="154" swimtime="00:00:40.53" resultid="5696" heatid="4793" lane="3" />
                <RESULT eventid="4425" points="165" swimtime="00:00:39.59" resultid="5730" heatid="4804" lane="6" />
                <RESULT eventid="4429" points="134" swimtime="00:00:43.14" resultid="5748" heatid="4853" lane="3" />
                <RESULT eventid="5807" points="121" swimtime="00:00:50.43" resultid="10124" heatid="6037" lane="3" />
                <RESULT eventid="5810" points="192" swimtime="00:00:34.94" resultid="10237" heatid="6021" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Mendes Costa" birthdate="2014-04-03" gender="F" nation="BRA" license="378341" swrid="5603873" athleteid="1729" externalid="378341" level="MRGA">
              <RESULTS>
                <RESULT eventid="1061" status="DNS" swimtime="00:00:00.00" resultid="1730" heatid="4654" lane="1" entrytime="00:00:54.62" entrycourse="SCM" />
                <RESULT eventid="1189" status="DNS" swimtime="00:00:00.00" resultid="1731" heatid="4935" lane="2" />
                <RESULT eventid="1298" status="DNS" swimtime="00:00:00.00" resultid="1732" heatid="5028" lane="6" entrytime="00:00:58.27" entrycourse="SCM" />
                <RESULT eventid="1311" status="DNS" swimtime="00:00:00.00" resultid="1733" heatid="5078" lane="4" entrytime="00:00:45.47" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Andrade Silva" birthdate="2016-03-15" gender="M" nation="BRA" license="414852" swrid="5755349" athleteid="1793" externalid="414852" level="MRGA">
              <RESULTS>
                <RESULT eventid="1201" points="89" swimtime="00:00:49.34" resultid="1794" heatid="4941" lane="3" entrytime="00:00:54.94" entrycourse="SCM" />
                <RESULT eventid="1225" points="76" swimtime="00:00:58.70" resultid="1795" heatid="4961" lane="3" entrytime="00:01:05.12" entrycourse="SCM" />
                <RESULT eventid="1261" points="111" swimtime="00:00:41.92" resultid="1796" heatid="4991" lane="3" entrytime="00:00:42.08" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Catarina" lastname="Wendt Jesus" birthdate="2013-07-09" gender="F" nation="BRA" license="393778" swrid="5641780" athleteid="1675" externalid="393778" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="306" swimtime="00:00:36.17" resultid="1676" heatid="4676" lane="3" entrytime="00:00:36.23" entrycourse="SCM" />
                <RESULT eventid="1077" points="288" swimtime="00:00:38.21" resultid="1677" heatid="4728" lane="5" entrytime="00:00:38.08" entrycourse="SCM" />
                <RESULT eventid="1179" points="344" swimtime="00:03:11.98" resultid="1678" heatid="4923" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.64" />
                    <SPLIT distance="100" swimtime="00:01:31.58" />
                    <SPLIT distance="150" swimtime="00:02:21.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="371" swimtime="00:01:09.92" resultid="1679" heatid="4938" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="322" swimtime="00:00:33.44" resultid="1680" heatid="5103" lane="6" entrytime="00:00:31.35" entrycourse="SCM" />
                <RESULT comment="SW 7.5 - Executou uma pernada de borboleta durante o nado.  (Horário: 8:38)" eventid="1301" status="DSQ" swimtime="00:00:41.77" resultid="1681" heatid="5051" lane="5" entrytime="00:00:40.83" entrycourse="SCM" />
                <RESULT eventid="4411" points="349" swimtime="00:00:34.60" resultid="5608" heatid="4679" lane="2" />
                <RESULT eventid="4413" points="362" swimtime="00:00:34.20" resultid="5633" heatid="4690" lane="4" />
                <RESULT eventid="4417" points="297" swimtime="00:00:37.83" resultid="5650" heatid="4730" lane="1" />
                <RESULT eventid="4419" points="335" swimtime="00:00:36.34" resultid="5677" heatid="4741" lane="4" />
                <RESULT eventid="5804" points="395" swimtime="00:00:31.24" resultid="10050" heatid="6053" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Casavechia Carraro" birthdate="2009-07-28" gender="M" nation="BRA" license="368150" swrid="5384752" athleteid="1418" externalid="368150" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="530" swimtime="00:00:26.86" resultid="1419" heatid="4782" lane="4" />
                <RESULT eventid="1105" points="273" swimtime="00:00:34.07" resultid="1420" heatid="4846" lane="6" />
                <RESULT eventid="1237" points="578" swimtime="00:00:57.33" resultid="1421" heatid="4977" lane="4" entrytime="00:00:58.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="642" swimtime="00:00:51.96" resultid="1422" heatid="5018" lane="4" entrytime="00:00:52.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="406" swimtime="00:00:27.21" resultid="1423" heatid="5226" lane="2" entrytime="00:00:24.99" entrycourse="SCM" />
                <RESULT eventid="1329" points="370" swimtime="00:00:34.74" resultid="1424" heatid="5160" lane="1" />
                <RESULT eventid="4423" points="415" swimtime="00:00:29.14" resultid="5716" heatid="4801" lane="1" />
                <RESULT eventid="4425" points="574" swimtime="00:00:26.16" resultid="5740" heatid="4808" lane="4" />
                <RESULT eventid="4429" points="328" swimtime="00:00:32.04" resultid="5766" heatid="4861" lane="1" />
                <RESULT eventid="4431" points="406" swimtime="00:00:29.85" resultid="5789" heatid="4868" lane="4" />
                <RESULT eventid="5807" points="411" swimtime="00:00:33.54" resultid="10143" heatid="6045" lane="1" />
                <RESULT eventid="5810" points="542" swimtime="00:00:24.72" resultid="10257" heatid="6029" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heitor" lastname="Bello Paula" birthdate="2015-06-14" gender="M" nation="BRA" license="393776" swrid="5507529" athleteid="1668" externalid="393776" level="MRGA">
              <RESULTS>
                <RESULT eventid="1089" points="72" swimtime="00:00:52.08" resultid="1669" heatid="4758" lane="1" entrytime="00:01:02.80" entrycourse="SCM" />
                <RESULT eventid="1102" points="87" swimtime="00:00:49.78" resultid="1670" heatid="4820" lane="1" entrytime="00:00:46.58" entrycourse="SCM" />
                <RESULT eventid="1213" points="93" swimtime="00:02:01.91" resultid="1671" heatid="4957" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="97" swimtime="00:01:37.57" resultid="1672" heatid="5013" lane="4" entrytime="00:01:37.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="110" swimtime="00:00:42.01" resultid="1673" heatid="5193" lane="5" entrytime="00:00:43.87" entrycourse="SCM" />
                <RESULT eventid="1326" points="84" swimtime="00:00:56.87" resultid="1674" heatid="5133" lane="6" entrytime="00:01:00.40" entrycourse="SCM" />
                <RESULT eventid="4427" points="82" swimtime="00:00:50.78" resultid="9030" heatid="9007" lane="6" />
                <RESULT eventid="4445" points="82" swimtime="00:00:57.23" resultid="10112" heatid="6033" lane="2" />
                <RESULT eventid="4451" points="120" swimtime="00:00:40.80" resultid="10225" heatid="6017" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Arthur Da Silva Ortiz" birthdate="2015-04-20" gender="M" nation="BRA" license="399733" swrid="5676285" athleteid="1696" externalid="399733" level="MRGA">
              <RESULTS>
                <RESULT eventid="1089" points="95" swimtime="00:00:47.53" resultid="1697" heatid="4759" lane="5" entrytime="00:00:48.66" entrycourse="SCM" />
                <RESULT eventid="1102" points="99" swimtime="00:00:47.65" resultid="1698" heatid="4819" lane="3" entrytime="00:00:51.54" entrycourse="SCM" />
                <RESULT eventid="1213" points="126" swimtime="00:01:50.06" resultid="1699" heatid="4956" lane="5" />
                <RESULT eventid="1237" points="69" swimtime="00:01:56.30" resultid="1700" heatid="4975" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="134" swimtime="00:00:39.34" resultid="1701" heatid="5193" lane="3" entrytime="00:00:41.36" entrycourse="SCM" />
                <RESULT eventid="1326" points="129" swimtime="00:00:49.28" resultid="1702" heatid="5134" lane="6" entrytime="00:00:52.04" entrycourse="SCM" />
                <RESULT eventid="4421" points="94" swimtime="00:00:47.78" resultid="9023" heatid="9005" lane="5" />
                <RESULT eventid="4427" points="96" swimtime="00:00:48.19" resultid="9029" heatid="9007" lane="5" />
                <RESULT eventid="4445" points="135" swimtime="00:00:48.59" resultid="10111" heatid="6033" lane="1" />
                <RESULT eventid="4451" points="138" swimtime="00:00:39.01" resultid="10223" heatid="6017" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Felipe Sakaguti" birthdate="2007-06-22" gender="M" nation="BRA" license="407187" swrid="5688778" athleteid="1750" externalid="407187" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="44" swimtime="00:01:01.28" resultid="1751" heatid="4783" lane="4" />
                <RESULT eventid="1105" points="93" swimtime="00:00:48.75" resultid="1752" heatid="4847" lane="1" entrytime="00:00:55.25" entrycourse="SCM" />
                <RESULT eventid="1273" points="106" swimtime="00:01:34.46" resultid="1753" heatid="5013" lane="3" entrytime="00:01:33.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="110" swimtime="00:00:42.03" resultid="1754" heatid="5219" lane="2" entrytime="00:00:42.66" entrycourse="SCM" />
                <RESULT comment="SW 7.5 - Executou uma pernada de borboleta durante o nado.  (Horário: 10:44)" eventid="1329" status="DSQ" swimtime="00:01:05.51" resultid="1755" heatid="5158" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Passafaro" birthdate="2009-02-01" gender="F" nation="BRA" license="370673" swrid="5603885" athleteid="1523" externalid="370673" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" status="DNS" swimtime="00:00:00.00" resultid="1524" heatid="4677" lane="2" entrytime="00:00:33.10" entrycourse="SCM" />
                <RESULT eventid="1077" status="DNS" swimtime="00:00:00.00" resultid="1525" heatid="4727" lane="3" entrytime="00:00:40.02" entrycourse="SCM" />
                <RESULT eventid="1153" status="DNS" swimtime="00:00:00.00" resultid="1526" heatid="4903" lane="4" entrytime="00:01:22.00" entrycourse="SCM" />
                <RESULT eventid="1189" status="DNS" swimtime="00:00:00.00" resultid="1527" heatid="4934" lane="4" entrytime="00:01:09.60" entrycourse="SCM" />
                <RESULT eventid="1314" status="DNS" swimtime="00:00:00.00" resultid="1528" heatid="5103" lane="5" entrytime="00:00:30.77" entrycourse="SCM" />
                <RESULT eventid="1301" status="DNS" swimtime="00:00:00.00" resultid="1529" heatid="5046" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Batista Sanchez" birthdate="2009-05-22" gender="M" nation="BRA" license="370668" swrid="5255779" athleteid="1439" externalid="370668" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="339" swimtime="00:00:31.19" resultid="1440" heatid="4789" lane="1" entrytime="00:00:34.73" entrycourse="SCM" />
                <RESULT eventid="1105" points="226" swimtime="00:00:36.29" resultid="1441" heatid="4843" lane="4" />
                <RESULT eventid="1213" points="389" swimtime="00:01:15.68" resultid="1442" heatid="4959" lane="5" entrytime="00:01:11.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="385" swimtime="00:02:45.14" resultid="1443" heatid="4995" lane="4" entrytime="00:02:41.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.63" />
                    <SPLIT distance="100" swimtime="00:01:19.89" />
                    <SPLIT distance="150" swimtime="00:02:02.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="345" swimtime="00:00:28.74" resultid="1444" heatid="5218" lane="2" />
                <RESULT eventid="1329" points="353" swimtime="00:00:35.28" resultid="1445" heatid="5165" lane="6" entrytime="00:00:34.30" entrycourse="SCM" />
                <RESULT eventid="4423" points="332" swimtime="00:00:31.38" resultid="5719" heatid="4801" lane="4" />
                <RESULT eventid="4429" points="201" swimtime="00:00:37.72" resultid="5769" heatid="4861" lane="4" />
                <RESULT eventid="5807" points="388" swimtime="00:00:34.18" resultid="10145" heatid="6045" lane="3" />
                <RESULT eventid="5810" points="342" swimtime="00:00:28.82" resultid="10259" heatid="6029" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lavinia" lastname="Bossoni" birthdate="2013-11-03" gender="F" nation="BRA" license="377260" swrid="5343093" athleteid="1565" externalid="377260" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="122" swimtime="00:00:49.14" resultid="1566" heatid="4675" lane="1" entrytime="00:00:46.76" entrycourse="SCM" />
                <RESULT eventid="1077" points="182" swimtime="00:00:44.54" resultid="1567" heatid="4726" lane="2" entrytime="00:00:43.59" entrycourse="SCM" />
                <RESULT eventid="1129" points="201" swimtime="00:01:46.35" resultid="1568" heatid="4889" lane="2" entrytime="00:01:46.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="203" swimtime="00:03:07.60" resultid="1569" heatid="4896" lane="2" entrytime="00:03:19.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.28" />
                    <SPLIT distance="100" swimtime="00:01:35.19" />
                    <SPLIT distance="150" swimtime="00:02:22.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="190" swimtime="00:00:39.86" resultid="1570" heatid="5099" lane="1" entrytime="00:00:39.07" entrycourse="SCM" />
                <RESULT eventid="1301" points="180" swimtime="00:00:50.19" resultid="1571" heatid="5049" lane="4" entrytime="00:00:51.39" entrycourse="SCM" />
                <RESULT eventid="4417" points="195" swimtime="00:00:43.53" resultid="5655" heatid="4730" lane="6" />
                <RESULT eventid="5801" points="180" swimtime="00:00:50.24" resultid="10013" heatid="6067" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathan" lastname="Novak Pinho" birthdate="2012-11-14" gender="M" nation="BRA" license="378199" swrid="5603879" athleteid="1593" externalid="378199" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="202" swimtime="00:00:37.04" resultid="1594" heatid="4785" lane="2" />
                <RESULT eventid="1105" points="186" swimtime="00:00:38.68" resultid="1595" heatid="4848" lane="4" entrytime="00:00:43.19" entrycourse="SCM" />
                <RESULT eventid="1288" points="235" swimtime="00:00:32.66" resultid="1596" heatid="5221" lane="6" entrytime="00:00:34.04" entrycourse="SCM" />
                <RESULT eventid="1329" points="112" swimtime="00:00:51.70" resultid="1597" heatid="5161" lane="3" />
                <RESULT eventid="4429" points="179" swimtime="00:00:39.23" resultid="5755" heatid="4855" lane="5" />
                <RESULT eventid="5810" points="224" swimtime="00:00:33.16" resultid="10245" heatid="6023" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Siqueira Almeida" birthdate="2016-06-21" gender="F" nation="BRA" license="414848" swrid="5755360" athleteid="1768" externalid="414848" level="MRGA">
              <RESULTS>
                <RESULT eventid="1117" points="110" swimtime="00:00:52.59" resultid="1769" heatid="4873" lane="3" entrytime="00:00:54.09" entrycourse="SCM" />
                <RESULT eventid="1141" points="75" swimtime="00:01:07.24" resultid="1770" heatid="4892" lane="3" entrytime="00:01:10.77" entrycourse="SCM" />
                <RESULT eventid="1177" points="64" swimtime="00:00:57.14" resultid="1771" heatid="4919" lane="3" entrytime="00:00:56.36" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Biason Santana" birthdate="2009-01-21" gender="M" nation="BRA" license="366969" swrid="5317765" athleteid="1537" externalid="366969" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="1538" heatid="4791" lane="5" entrytime="00:00:27.47" entrycourse="SCM" />
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="1539" heatid="4844" lane="2" />
                <RESULT eventid="1237" status="DNS" swimtime="00:00:00.00" resultid="1540" heatid="4975" lane="3" entrytime="00:01:02.60" entrycourse="SCM" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="1541" heatid="5017" lane="3" entrytime="00:00:58.82" entrycourse="SCM" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="1542" heatid="5225" lane="1" entrytime="00:00:27.49" entrycourse="SCM" />
                <RESULT eventid="1329" status="DNS" swimtime="00:00:00.00" resultid="1543" heatid="5158" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Dos Reis Monteiro" birthdate="2014-08-05" gender="M" nation="BRA" license="392095" swrid="5697226" athleteid="1619" externalid="392095" level="MRGA">
              <RESULTS>
                <RESULT eventid="1089" points="214" swimtime="00:00:36.31" resultid="1620" heatid="4759" lane="3" entrytime="00:00:37.00" entrycourse="SCM" />
                <RESULT eventid="1102" points="144" swimtime="00:00:42.18" resultid="1621" heatid="4820" lane="2" entrytime="00:00:45.97" entrycourse="SCM" />
                <RESULT eventid="1213" points="196" swimtime="00:01:35.13" resultid="1622" heatid="4955" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="213" swimtime="00:01:15.01" resultid="1623" heatid="5015" lane="2" entrytime="00:01:15.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="205" swimtime="00:00:34.16" resultid="1624" heatid="5194" lane="3" entrytime="00:00:32.22" entrycourse="SCM" />
                <RESULT eventid="1326" points="190" swimtime="00:00:43.36" resultid="1625" heatid="5134" lane="3" entrytime="00:00:40.93" entrycourse="SCM" />
                <RESULT eventid="4421" points="227" swimtime="00:00:35.64" resultid="9025" heatid="9006" lane="4" />
                <RESULT eventid="4427" points="152" swimtime="00:00:41.41" resultid="9031" heatid="9008" lane="4" />
                <RESULT eventid="4445" points="207" swimtime="00:00:42.11" resultid="10116" heatid="6035" lane="1" />
                <RESULT eventid="4451" points="216" swimtime="00:00:33.55" resultid="10229" heatid="6019" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carina" lastname="Costa Profeta" birthdate="2008-03-20" gender="F" nation="BRA" license="366964" swrid="5591584" athleteid="1509" externalid="366964" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="457" swimtime="00:00:31.63" resultid="1510" heatid="4672" lane="2" />
                <RESULT eventid="1077" points="288" swimtime="00:00:38.22" resultid="1511" heatid="4724" lane="2" />
                <RESULT eventid="1129" points="482" swimtime="00:01:19.51" resultid="1512" heatid="4890" lane="3" entrytime="00:01:19.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="393" swimtime="00:01:08.55" resultid="1513" heatid="4939" lane="2" entrytime="00:01:05.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="223" swimtime="00:00:37.77" resultid="1514" heatid="5103" lane="1" entrytime="00:00:30.78" entrycourse="SCM" />
                <RESULT eventid="1301" points="443" swimtime="00:00:37.20" resultid="1515" heatid="5051" lane="3" entrytime="00:00:35.68" entrycourse="SCM" />
                <RESULT eventid="4411" points="398" swimtime="00:00:33.12" resultid="5630" heatid="4689" lane="1" />
                <RESULT eventid="4413" points="465" swimtime="00:00:31.45" resultid="5647" heatid="4695" lane="4" />
                <RESULT eventid="4417" points="279" swimtime="00:00:38.64" resultid="5673" heatid="4740" lane="1" />
                <RESULT eventid="4419" points="338" swimtime="00:00:36.24" resultid="5691" heatid="4746" lane="4" />
                <RESULT eventid="5801" points="425" swimtime="00:00:37.72" resultid="10036" heatid="6077" lane="1" />
                <RESULT eventid="5804" points="390" swimtime="00:00:31.36" resultid="10076" heatid="6063" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Meneghetti Vidal" birthdate="2015-06-12" gender="M" nation="BRA" license="414851" swrid="5757894" athleteid="1786" externalid="414851" level="MRGA">
              <RESULTS>
                <RESULT eventid="1089" points="62" swimtime="00:00:54.77" resultid="1787" heatid="4758" lane="5" entrytime="00:00:58.49" entrycourse="SCM" />
                <RESULT eventid="1102" points="69" swimtime="00:00:53.84" resultid="1788" heatid="4819" lane="2" entrytime="00:00:57.71" entrycourse="SCM" />
                <RESULT eventid="1237" points="51" swimtime="00:02:08.03" resultid="1789" heatid="4975" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="104" swimtime="00:01:35.24" resultid="1790" heatid="5012" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="103" swimtime="00:00:43.00" resultid="1791" heatid="5193" lane="6" entrytime="00:00:44.86" entrycourse="SCM" />
                <RESULT eventid="1326" points="58" swimtime="00:01:04.32" resultid="1792" heatid="5132" lane="4" entrytime="00:01:04.01" entrycourse="SCM" />
                <RESULT eventid="4445" points="63" swimtime="00:01:02.38" resultid="10115" heatid="6033" lane="5" />
                <RESULT eventid="4451" points="106" swimtime="00:00:42.56" resultid="10226" heatid="6017" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabrielle" lastname="Borba" birthdate="2014-06-15" gender="F" nation="BRA" license="385705" swrid="5323267" athleteid="1612" externalid="385705" level="MRGA">
              <RESULTS>
                <RESULT eventid="1061" points="118" swimtime="00:00:49.57" resultid="1613" heatid="4653" lane="5" />
                <RESULT eventid="1074" points="119" swimtime="00:00:51.31" resultid="1614" heatid="4705" lane="6" entrytime="00:00:53.78" entrycourse="SCM" />
                <RESULT eventid="1129" points="147" swimtime="00:01:57.90" resultid="1615" heatid="4889" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="150" swimtime="00:01:34.48" resultid="1616" heatid="4935" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="131" swimtime="00:00:55.86" resultid="1617" heatid="5028" lane="2" entrytime="00:00:54.15" entrycourse="SCM" />
                <RESULT eventid="1311" points="161" swimtime="00:00:42.10" resultid="1618" heatid="5079" lane="1" entrytime="00:00:41.54" entrycourse="SCM" />
                <RESULT eventid="4409" points="132" swimtime="00:00:47.88" resultid="9020" heatid="9002" lane="6" />
                <RESULT eventid="4433" points="139" swimtime="00:00:54.68" resultid="10007" heatid="6065" lane="3" />
                <RESULT eventid="4439" points="172" swimtime="00:00:41.21" resultid="10047" heatid="6051" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juan" lastname="Bernardo Padua" birthdate="2013-07-15" gender="M" nation="BRA" license="392108" swrid="5305422" athleteid="1640" externalid="392108" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="179" swimtime="00:00:38.55" resultid="1641" heatid="4787" lane="3" entrytime="00:00:38.33" entrycourse="SCM" />
                <RESULT eventid="1105" points="115" swimtime="00:00:45.37" resultid="1642" heatid="4848" lane="3" entrytime="00:00:42.43" entrycourse="SCM" />
                <RESULT eventid="1213" points="179" swimtime="00:01:37.93" resultid="1643" heatid="4958" lane="1" entrytime="00:01:38.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="176" swimtime="00:03:34.40" resultid="1644" heatid="4995" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.24" />
                    <SPLIT distance="100" swimtime="00:01:45.43" />
                    <SPLIT distance="150" swimtime="00:02:42.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="193" swimtime="00:00:34.88" resultid="1645" heatid="5220" lane="5" entrytime="00:00:35.98" entrycourse="SCM" />
                <RESULT eventid="1329" points="177" swimtime="00:00:44.39" resultid="1646" heatid="5163" lane="2" entrytime="00:00:44.56" entrycourse="SCM" />
                <RESULT eventid="4423" points="165" swimtime="00:00:39.60" resultid="5695" heatid="4793" lane="2" />
                <RESULT eventid="4425" points="165" swimtime="00:00:39.62" resultid="5729" heatid="4804" lane="5" />
                <RESULT eventid="4429" points="151" swimtime="00:00:41.46" resultid="5749" heatid="4853" lane="4" />
                <RESULT eventid="4431" points="148" swimtime="00:00:41.72" resultid="5778" heatid="4864" lane="5" />
                <RESULT eventid="5807" points="191" swimtime="00:00:43.32" resultid="10122" heatid="6037" lane="1" />
                <RESULT eventid="5810" points="196" swimtime="00:00:34.66" resultid="10236" heatid="6021" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Pavão" birthdate="2012-04-04" gender="F" nation="BRA" license="377259" swrid="5603888" athleteid="1558" externalid="377259" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="234" swimtime="00:00:39.55" resultid="1559" heatid="4676" lane="6" entrytime="00:00:40.84" entrycourse="SCM" />
                <RESULT eventid="1077" points="263" swimtime="00:00:39.37" resultid="1560" heatid="4727" lane="2" entrytime="00:00:40.95" entrycourse="SCM" />
                <RESULT eventid="1119" points="305" swimtime="00:02:56.63" resultid="1561" heatid="4878" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.15" />
                    <SPLIT distance="100" swimtime="00:01:27.06" />
                    <SPLIT distance="150" swimtime="00:02:12.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="291" swimtime="00:01:22.83" resultid="1562" heatid="4917" lane="5" entrytime="00:01:23.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="307" swimtime="00:00:33.98" resultid="1563" heatid="5101" lane="6" entrytime="00:00:34.35" entrycourse="SCM" />
                <RESULT eventid="1301" points="252" swimtime="00:00:44.90" resultid="1564" heatid="5050" lane="5" entrytime="00:00:47.46" entrycourse="SCM" />
                <RESULT eventid="4411" points="240" swimtime="00:00:39.21" resultid="5616" heatid="4681" lane="4" />
                <RESULT eventid="4413" points="241" swimtime="00:00:39.15" resultid="5638" heatid="4691" lane="6" />
                <RESULT eventid="4417" points="284" swimtime="00:00:38.37" resultid="5658" heatid="4732" lane="3" />
                <RESULT eventid="4419" points="280" swimtime="00:00:38.59" resultid="5682" heatid="4742" lane="6" />
                <RESULT eventid="5801" points="241" swimtime="00:00:45.53" resultid="10021" heatid="6069" lane="5" />
                <RESULT eventid="5804" points="313" swimtime="00:00:33.77" resultid="10058" heatid="6055" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Ayres" birthdate="2012-05-05" gender="M" nation="BRA" license="378035" swrid="5208079" athleteid="1586" externalid="378035" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="285" swimtime="00:00:33.02" resultid="1587" heatid="4789" lane="3" entrytime="00:00:32.81" entrycourse="SCM" />
                <RESULT eventid="1105" points="234" swimtime="00:00:35.87" resultid="1588" heatid="4850" lane="5" entrytime="00:00:34.60" entrycourse="SCM" />
                <RESULT eventid="1203" points="261" swimtime="00:02:45.14" resultid="1589" heatid="4944" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                    <SPLIT distance="100" swimtime="00:01:22.33" />
                    <SPLIT distance="150" swimtime="00:02:05.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1237" points="256" swimtime="00:01:15.22" resultid="1590" heatid="4976" lane="4" entrytime="00:01:14.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="269" swimtime="00:00:31.20" resultid="1591" heatid="5223" lane="6" entrytime="00:00:30.93" entrycourse="SCM" />
                <RESULT eventid="1329" points="241" swimtime="00:00:40.08" resultid="1592" heatid="5164" lane="6" entrytime="00:00:41.70" entrycourse="SCM" />
                <RESULT eventid="4423" points="290" swimtime="00:00:32.85" resultid="5700" heatid="4795" lane="2" />
                <RESULT eventid="4425" points="298" swimtime="00:00:32.53" resultid="5732" heatid="4805" lane="5" />
                <RESULT eventid="4429" points="249" swimtime="00:00:35.10" resultid="5751" heatid="4855" lane="1" />
                <RESULT eventid="4431" points="275" swimtime="00:00:33.97" resultid="5780" heatid="4865" lane="4" />
                <RESULT eventid="5807" points="240" swimtime="00:00:40.12" resultid="10127" heatid="6039" lane="1" />
                <RESULT eventid="5810" points="301" swimtime="00:00:30.08" resultid="10240" heatid="6023" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Schuch Pimpao" birthdate="2010-05-17" gender="M" nation="BRA" license="355586" swrid="5588908" athleteid="1467" externalid="355586" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="290" swimtime="00:00:32.85" resultid="1468" heatid="4783" lane="3" />
                <RESULT eventid="1105" points="249" swimtime="00:00:35.11" resultid="1469" heatid="4850" lane="4" entrytime="00:00:31.29" entrycourse="SCM" />
                <RESULT eventid="1203" points="370" swimtime="00:02:27.05" resultid="1470" heatid="4945" lane="4" entrytime="00:02:28.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                    <SPLIT distance="100" swimtime="00:01:10.98" />
                    <SPLIT distance="150" swimtime="00:01:49.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="357" swimtime="00:01:08.11" resultid="1471" heatid="4989" lane="2" entrytime="00:01:08.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="262" swimtime="00:00:31.49" resultid="1472" heatid="5217" lane="2" />
                <RESULT eventid="1329" points="270" swimtime="00:00:38.56" resultid="1473" heatid="5159" lane="4" />
                <RESULT eventid="4423" points="265" swimtime="00:00:33.86" resultid="5714" heatid="4799" lane="2" />
                <RESULT eventid="4425" points="301" swimtime="00:00:32.44" resultid="5738" heatid="4807" lane="5" />
                <RESULT eventid="4429" points="212" swimtime="00:00:37.06" resultid="5763" heatid="4859" lane="1" />
                <RESULT eventid="4431" points="341" swimtime="00:00:31.62" resultid="5786" heatid="4867" lane="4" />
                <RESULT eventid="5807" points="286" swimtime="00:00:37.86" resultid="10141" heatid="6043" lane="2" />
                <RESULT eventid="5810" points="365" swimtime="00:00:28.20" resultid="10253" heatid="6027" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Pastre" birthdate="2014-03-10" gender="F" nation="BRA" license="403760" swrid="5684593" athleteid="1722" externalid="403760" level="MRGA">
              <RESULTS>
                <RESULT eventid="1061" points="171" swimtime="00:00:43.88" resultid="1723" heatid="4654" lane="2" entrytime="00:00:45.93" entrycourse="SCM" />
                <RESULT eventid="1074" points="228" swimtime="00:00:41.32" resultid="1724" heatid="4705" lane="3" entrytime="00:00:40.11" entrycourse="SCM" />
                <RESULT eventid="1165" points="196" swimtime="00:01:34.44" resultid="1725" heatid="4915" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="193" swimtime="00:01:26.95" resultid="1726" heatid="4936" lane="4" entrytime="00:01:46.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="139" swimtime="00:00:54.71" resultid="1727" heatid="5028" lane="1" entrytime="00:00:55.79" entrycourse="SCM" />
                <RESULT eventid="1311" points="189" swimtime="00:00:39.90" resultid="1728" heatid="5079" lane="4" entrytime="00:00:37.81" entrycourse="SCM" />
                <RESULT eventid="4415" points="250" swimtime="00:00:40.03" resultid="9013" heatid="9004" lane="4" />
                <RESULT eventid="4409" points="162" swimtime="00:00:44.65" resultid="9019" heatid="9002" lane="5" />
                <RESULT eventid="4433" points="150" swimtime="00:00:53.38" resultid="10006" heatid="6065" lane="2" />
                <RESULT eventid="4439" points="191" swimtime="00:00:39.81" resultid="10045" heatid="6051" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kauan" lastname="Gabriel Pereira" birthdate="2014-05-14" gender="M" nation="BRA" license="407181" swrid="5718625" athleteid="1743" externalid="407181" level="MRGA">
              <RESULTS>
                <RESULT eventid="1089" points="66" swimtime="00:00:53.78" resultid="1744" heatid="4758" lane="2" entrytime="00:00:58.30" entrycourse="SCM" />
                <RESULT eventid="1102" points="90" swimtime="00:00:49.32" resultid="1745" heatid="4819" lane="4" entrytime="00:00:51.63" entrycourse="SCM" />
                <RESULT eventid="1249" points="94" swimtime="00:01:46.00" resultid="1746" heatid="4987" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="107" swimtime="00:01:34.33" resultid="1747" heatid="5013" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="107" swimtime="00:00:42.46" resultid="1748" heatid="5193" lane="1" entrytime="00:00:44.61" entrycourse="SCM" />
                <RESULT eventid="1326" points="75" swimtime="00:00:59.00" resultid="1749" heatid="5132" lane="2" entrytime="00:01:32.58" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Mochiutti Carneiro" birthdate="2010-04-22" gender="F" nation="BRA" license="370670" swrid="5588817" athleteid="1481" externalid="370670" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="378" swimtime="00:00:33.69" resultid="1482" heatid="4677" lane="3" entrytime="00:00:31.98" entrycourse="SCM" />
                <RESULT eventid="1077" points="286" swimtime="00:00:38.31" resultid="1483" heatid="4723" lane="3" />
                <RESULT eventid="1143" points="432" swimtime="00:02:25.81" resultid="1484" heatid="4897" lane="3" entrytime="00:02:21.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                    <SPLIT distance="100" swimtime="00:01:10.24" />
                    <SPLIT distance="150" swimtime="00:01:48.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="437" swimtime="00:01:06.20" resultid="1485" heatid="4939" lane="3" entrytime="00:01:03.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="241" swimtime="00:00:36.80" resultid="1486" heatid="5103" lane="4" entrytime="00:00:29.36" entrycourse="SCM" />
                <RESULT eventid="1301" points="268" swimtime="00:00:43.99" resultid="1487" heatid="5046" lane="2" />
                <RESULT eventid="4411" points="388" swimtime="00:00:33.40" resultid="5624" heatid="4685" lane="2" />
                <RESULT eventid="4413" points="415" swimtime="00:00:32.66" resultid="5642" heatid="4693" lane="4" />
                <RESULT eventid="4417" points="312" swimtime="00:00:37.22" resultid="5668" heatid="4736" lane="3" />
                <RESULT eventid="4419" points="325" swimtime="00:00:36.69" resultid="5686" heatid="4744" lane="4" />
                <RESULT eventid="5801" points="287" swimtime="00:00:42.99" resultid="10028" heatid="6073" lane="2" />
                <RESULT eventid="5804" points="422" swimtime="00:00:30.57" resultid="10071" heatid="6059" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1115" points="297" swimtime="00:04:28.78" resultid="1803" heatid="5251" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.88" />
                    <SPLIT distance="100" swimtime="00:01:10.15" />
                    <SPLIT distance="150" swimtime="00:01:40.66" />
                    <SPLIT distance="200" swimtime="00:02:26.89" />
                    <SPLIT distance="250" swimtime="00:03:02.94" />
                    <SPLIT distance="300" swimtime="00:03:34.68" />
                    <SPLIT distance="350" swimtime="00:04:01.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1696" number="1" />
                    <RELAYPOSITION athleteid="1530" number="2" />
                    <RELAYPOSITION athleteid="1467" number="3" />
                    <RELAYPOSITION athleteid="1640" number="4" />
                    <RELAYPOSITION athleteid="1619" number="5" />
                    <RELAYPOSITION athleteid="1586" number="6" />
                    <RELAYPOSITION athleteid="1405" number="7" />
                    <RELAYPOSITION athleteid="1418" number="8" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1339" points="305" swimtime="00:04:02.90" resultid="10109" heatid="5252" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.05" />
                    <SPLIT distance="100" swimtime="00:01:09.35" />
                    <SPLIT distance="150" swimtime="00:01:45.14" />
                    <SPLIT distance="200" swimtime="00:02:19.41" />
                    <SPLIT distance="250" swimtime="00:02:45.79" />
                    <SPLIT distance="300" swimtime="00:03:13.14" />
                    <SPLIT distance="350" swimtime="00:03:37.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1586" number="1" />
                    <RELAYPOSITION athleteid="1696" number="2" />
                    <RELAYPOSITION athleteid="1640" number="3" />
                    <RELAYPOSITION athleteid="1619" number="4" />
                    <RELAYPOSITION athleteid="1405" number="5" />
                    <RELAYPOSITION athleteid="1467" number="6" />
                    <RELAYPOSITION athleteid="1418" number="7" />
                    <RELAYPOSITION athleteid="1432" number="8" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="APAN MARINGÁ &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1115" points="227" status="EXH" swimtime="00:04:53.77" resultid="5795" heatid="5251" lane="5" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.60" />
                    <SPLIT distance="100" swimtime="00:01:25.44" />
                    <SPLIT distance="150" swimtime="00:02:05.26" />
                    <SPLIT distance="200" swimtime="00:02:34.19" />
                    <SPLIT distance="250" swimtime="00:03:12.08" />
                    <SPLIT distance="300" swimtime="00:03:51.88" />
                    <SPLIT distance="350" swimtime="00:04:26.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1626" number="1" />
                    <RELAYPOSITION athleteid="1682" number="2" />
                    <RELAYPOSITION athleteid="1654" number="3" />
                    <RELAYPOSITION athleteid="1572" number="4" />
                    <RELAYPOSITION athleteid="1453" number="5" />
                    <RELAYPOSITION athleteid="1460" number="6" />
                    <RELAYPOSITION athleteid="1439" number="7" />
                    <RELAYPOSITION athleteid="1405" number="8" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="APAN/MARINGÁ &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1339" points="266" status="EXH" swimtime="00:04:14.21" resultid="1804" heatid="5252" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="100" swimtime="00:01:07.70" />
                    <SPLIT distance="150" swimtime="00:01:47.27" />
                    <SPLIT distance="200" swimtime="00:02:21.50" />
                    <SPLIT distance="250" swimtime="00:02:51.45" />
                    <SPLIT distance="300" swimtime="00:03:21.29" />
                    <SPLIT distance="350" swimtime="00:03:48.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1460" number="1" />
                    <RELAYPOSITION athleteid="1682" number="2" />
                    <RELAYPOSITION athleteid="1668" number="3" />
                    <RELAYPOSITION athleteid="1654" number="4" />
                    <RELAYPOSITION athleteid="1453" number="5" />
                    <RELAYPOSITION athleteid="1572" number="6" />
                    <RELAYPOSITION athleteid="1439" number="7" />
                    <RELAYPOSITION athleteid="1530" number="8" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT comment="SW 10.12 - Os pés perderam contato com a plataforma de partida antes que o colega de equipe anterior tocasse a borda.  (Horário: 11:20)" eventid="1087" status="DSQ" swimtime="00:05:17.08" resultid="1801" heatid="5247" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.78" />
                    <SPLIT distance="100" swimtime="00:01:44.62" />
                    <SPLIT distance="150" swimtime="00:02:19.36" />
                    <SPLIT distance="200" swimtime="00:03:01.01" />
                    <SPLIT distance="250" swimtime="00:03:32.25" />
                    <SPLIT distance="300" swimtime="00:04:05.10" />
                    <SPLIT distance="350" swimtime="00:04:36.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1675" number="1" />
                    <RELAYPOSITION athleteid="1734" number="2" />
                    <RELAYPOSITION athleteid="1516" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="1598" number="4" status="DSQ" />
                    <RELAYPOSITION athleteid="1509" number="5" status="DSQ" />
                    <RELAYPOSITION athleteid="1481" number="6" status="DSQ" />
                    <RELAYPOSITION athleteid="1488" number="7" status="DSQ" />
                    <RELAYPOSITION athleteid="1722" number="8" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1324" points="305" swimtime="00:04:34.78" resultid="1802" heatid="5249" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                    <SPLIT distance="100" swimtime="00:01:18.82" />
                    <SPLIT distance="150" swimtime="00:01:58.74" />
                    <SPLIT distance="200" swimtime="00:02:30.81" />
                    <SPLIT distance="250" swimtime="00:03:00.41" />
                    <SPLIT distance="300" swimtime="00:03:31.35" />
                    <SPLIT distance="350" swimtime="00:04:04.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1558" number="1" />
                    <RELAYPOSITION athleteid="1772" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1722" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1488" number="4" reactiontime="0" />
                    <RELAYPOSITION athleteid="1481" number="5" reactiontime="0" />
                    <RELAYPOSITION athleteid="1675" number="6" reactiontime="0" />
                    <RELAYPOSITION athleteid="1516" number="7" reactiontime="0" />
                    <RELAYPOSITION athleteid="1509" number="8" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="2539" nation="BRA" region="PR" clubid="2131" swrid="93771" name="Círculo Militar Do Paraná" shortname="Círculo Militar">
          <ATHLETES>
            <ATHLETE firstname="Vicente" lastname="Bileski" birthdate="2011-06-29" gender="M" nation="BRA" license="406950" swrid="5717248" athleteid="2167" externalid="406950" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="248" swimtime="00:00:34.59" resultid="2168" heatid="4772" lane="3" />
                <RESULT eventid="1105" points="174" swimtime="00:00:39.58" resultid="2169" heatid="4831" lane="1" />
                <RESULT eventid="1237" points="226" swimtime="00:01:18.41" resultid="2170" heatid="4971" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="275" swimtime="00:01:08.92" resultid="2171" heatid="4998" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente., Na volta dos 25m." eventid="1329" status="DSQ" swimtime="00:00:43.39" resultid="2173" heatid="5150" lane="5" entrytime="00:00:47.91" entrycourse="SCM" />
                <RESULT eventid="10332" points="259" swimtime="00:00:31.62" resultid="10398" heatid="10350" lane="2" entrytime="00:00:37.67" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Manocchio" birthdate="2011-07-28" gender="M" nation="BRA" license="384916" swrid="5588573" athleteid="2160" externalid="384916" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="247" swimtime="00:00:34.65" resultid="2161" heatid="4777" lane="6" entrytime="00:00:37.33" entrycourse="SCM" />
                <RESULT eventid="1105" points="229" swimtime="00:00:36.10" resultid="2162" heatid="4824" lane="1" />
                <RESULT eventid="1227" points="398" swimtime="00:02:15.04" resultid="2163" heatid="4964" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                    <SPLIT distance="100" swimtime="00:01:05.18" />
                    <SPLIT distance="150" swimtime="00:01:40.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="375" swimtime="00:01:02.16" resultid="2164" heatid="5008" lane="1" entrytime="00:01:05.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="236" swimtime="00:00:40.32" resultid="2166" heatid="5144" lane="5" />
                <RESULT eventid="10332" points="355" swimtime="00:00:28.46" resultid="10397" heatid="10356" lane="4" entrytime="00:00:29.60" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Maria Romanelli" birthdate="2011-04-18" gender="F" nation="BRA" license="378335" swrid="5588803" athleteid="2153" externalid="378335" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="242" swimtime="00:00:39.08" resultid="2154" heatid="4665" lane="5" />
                <RESULT eventid="1077" points="249" swimtime="00:00:40.12" resultid="2155" heatid="4719" lane="6" entrytime="00:00:40.11" entrycourse="SCM" />
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="2156" heatid="4908" lane="3" />
                <RESULT eventid="1189" status="DNS" swimtime="00:00:00.00" resultid="2157" heatid="4931" lane="4" entrytime="00:01:10.00" entrycourse="SCM" />
                <RESULT eventid="1314" points="363" swimtime="00:00:32.14" resultid="2158" heatid="5093" lane="1" entrytime="00:00:32.35" entrycourse="SCM" />
                <RESULT eventid="1301" points="249" swimtime="00:00:45.08" resultid="2159" heatid="5041" lane="1" entrytime="00:00:47.46" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Vieira De Macedo Brasil" birthdate="2009-12-19" gender="F" nation="BRA" license="344143" swrid="5622311" athleteid="2139" externalid="344143" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="246" swimtime="00:00:38.86" resultid="2140" heatid="4661" lane="4" />
                <RESULT eventid="1077" points="217" swimtime="00:00:41.96" resultid="2141" heatid="4712" lane="5" />
                <RESULT eventid="1179" points="304" swimtime="00:03:20.01" resultid="2142" heatid="4920" lane="2" />
                <RESULT eventid="1143" points="400" swimtime="00:02:29.64" resultid="2143" heatid="4893" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="383" swimtime="00:00:31.57" resultid="2144" heatid="5093" lane="2" entrytime="00:00:32.11" entrycourse="SCM" />
                <RESULT eventid="1301" points="323" swimtime="00:00:41.34" resultid="2145" heatid="5042" lane="7" entrytime="00:00:42.51" entrycourse="SCM" />
                <RESULT eventid="5801" points="336" swimtime="00:00:40.79" resultid="10544" heatid="6074" lane="5" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernando" lastname="Jun Melo Ogima" birthdate="2006-07-05" gender="M" nation="BRA" license="378332" swrid="5622284" athleteid="2146" externalid="378332" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="341" swimtime="00:00:31.13" resultid="2147" heatid="4780" lane="6" entrytime="00:00:30.48" entrycourse="SCM" />
                <RESULT eventid="1105" points="294" swimtime="00:00:33.23" resultid="2148" heatid="4840" lane="2" entrytime="00:00:33.73" entrycourse="SCM" />
                <RESULT eventid="1237" points="258" swimtime="00:01:14.96" resultid="2149" heatid="4969" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="366" swimtime="00:01:02.63" resultid="2150" heatid="4997" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="309" swimtime="00:00:36.87" resultid="2152" heatid="5155" lane="8" entrytime="00:00:35.92" entrycourse="SCM" />
                <RESULT eventid="10332" points="376" swimtime="00:00:27.92" resultid="10396" heatid="10359" lane="8" entrytime="00:00:27.54" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathan" lastname="Torres Oliveira" birthdate="2008-04-10" gender="M" nation="BRA" license="400274" swrid="5653303" athleteid="2132" externalid="400274" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="391" swimtime="00:00:29.74" resultid="2133" heatid="4766" lane="6" />
                <RESULT eventid="1105" points="278" swimtime="00:00:33.85" resultid="2134" heatid="4839" lane="6" entrytime="00:00:36.71" entrycourse="SCM" />
                <RESULT eventid="1249" points="248" swimtime="00:01:16.86" resultid="2135" heatid="4983" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="399" swimtime="00:01:00.89" resultid="2136" heatid="5007" lane="5" entrytime="00:01:07.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="311" swimtime="00:00:36.82" resultid="2138" heatid="5154" lane="5" entrytime="00:00:37.39" entrycourse="SCM" />
                <RESULT eventid="10332" points="428" swimtime="00:00:26.75" resultid="10395" heatid="10357" lane="1" entrytime="00:00:29.24" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2864" nation="BRA" region="PR" clubid="1341" swrid="93756" name="Associacao De Pais E Amigos Da Natacao De Ponta Gr" shortname="Apan Ponta Grossa">
          <ATHLETES>
            <ATHLETE firstname="Ana" lastname="Clara Domingues" birthdate="2012-01-19" gender="F" nation="BRA" license="377291" swrid="5588599" athleteid="1370" externalid="377291" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="87" swimtime="00:00:54.90" resultid="1371" heatid="4659" lane="5" />
                <RESULT eventid="1077" points="186" swimtime="00:00:44.20" resultid="1372" heatid="4715" lane="5" entrytime="00:00:49.20" entrycourse="SCM" />
                <RESULT eventid="1165" points="178" swimtime="00:01:37.40" resultid="1373" heatid="4912" lane="5" entrytime="00:01:36.16" entrycourse="SCM" />
                <RESULT eventid="1189" points="239" swimtime="00:01:20.89" resultid="1374" heatid="4929" lane="4" entrytime="00:01:18.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="234" swimtime="00:00:37.18" resultid="1375" heatid="5084" lane="1" />
                <RESULT eventid="1301" points="88" swimtime="00:01:03.65" resultid="1376" heatid="5031" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolly" lastname="Victoria Souza" birthdate="2015-11-15" gender="F" nation="BRA" license="400091" swrid="5652902" athleteid="1391" externalid="400091" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="79" swimtime="00:00:56.63" resultid="1392" heatid="4646" lane="1" />
                <RESULT eventid="1074" points="116" swimtime="00:00:51.73" resultid="1393" heatid="4698" lane="1" entrytime="00:00:57.81" entrycourse="SCM" />
                <RESULT eventid="1129" points="146" swimtime="00:01:58.24" resultid="1394" heatid="4884" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="136" swimtime="00:00:55.16" resultid="1395" heatid="5024" lane="4" entrytime="00:00:55.66" entrycourse="SCM" />
                <RESULT eventid="1311" points="143" swimtime="00:00:43.83" resultid="1396" heatid="5073" lane="6" entrytime="00:00:44.61" entrycourse="SCM" />
                <RESULT eventid="4415" points="112" swimtime="00:00:52.34" resultid="5401" heatid="4706" lane="6" />
                <RESULT eventid="4433" points="136" swimtime="00:00:55.14" resultid="10084" heatid="5029" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Chi Kravchychyn" birthdate="2009-09-27" gender="M" nation="BRA" license="344268" swrid="5600134" athleteid="1342" externalid="344268" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="478" swimtime="00:00:27.81" resultid="1343" heatid="4781" lane="1" entrytime="00:00:28.33" entrycourse="SCM" />
                <RESULT eventid="1105" points="361" swimtime="00:00:31.05" resultid="1344" heatid="4840" lane="3" entrytime="00:00:31.60" entrycourse="SCM" />
                <RESULT eventid="1203" points="432" swimtime="00:02:19.69" resultid="1345" heatid="4942" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                    <SPLIT distance="100" swimtime="00:01:09.57" />
                    <SPLIT distance="150" swimtime="00:01:45.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="510" swimtime="00:02:04.37" resultid="1346" heatid="4962" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.45" />
                    <SPLIT distance="100" swimtime="00:00:59.86" />
                    <SPLIT distance="150" swimtime="00:01:32.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="487" swimtime="00:00:31.70" resultid="1348" heatid="5155" lane="3" entrytime="00:00:32.19" entrycourse="SCM" />
                <RESULT eventid="4423" points="445" swimtime="00:00:28.47" resultid="5549" heatid="4800" lane="3" />
                <RESULT eventid="4429" points="367" swimtime="00:00:30.87" resultid="5588" heatid="4860" lane="4" />
                <RESULT eventid="5807" points="482" swimtime="00:00:31.80" resultid="10294" heatid="6044" lane="3" />
                <RESULT eventid="10332" points="487" swimtime="00:00:25.62" resultid="10361" heatid="10348" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Miretzki" birthdate="2014-09-17" gender="F" nation="BRA" license="414996" swrid="5755341" athleteid="1397" externalid="414996" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="89" swimtime="00:00:54.47" resultid="1398" heatid="4645" lane="2" />
                <RESULT eventid="1074" points="126" swimtime="00:00:50.32" resultid="1399" heatid="4697" lane="1" />
                <RESULT eventid="1298" points="134" swimtime="00:00:55.35" resultid="1400" heatid="5020" lane="8" />
                <RESULT eventid="1311" points="216" swimtime="00:00:38.16" resultid="1401" heatid="5072" lane="7" />
                <RESULT eventid="4439" points="222" swimtime="00:00:37.84" resultid="10185" heatid="6050" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Fegert" birthdate="2009-04-13" gender="M" nation="BRA" license="353813" swrid="5622279" athleteid="1363" externalid="353813" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="479" swimtime="00:00:27.79" resultid="1364" heatid="4781" lane="6" entrytime="00:00:28.38" entrycourse="SCM" />
                <RESULT eventid="1105" points="342" swimtime="00:00:31.60" resultid="1365" heatid="4828" lane="2" />
                <RESULT eventid="1237" points="432" swimtime="00:01:03.20" resultid="1366" heatid="4974" lane="4" entrytime="00:01:02.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="433" swimtime="00:00:59.24" resultid="1367" heatid="5011" lane="1" entrytime="00:00:57.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="347" swimtime="00:00:35.50" resultid="1369" heatid="5147" lane="3" />
                <RESULT eventid="4423" points="474" swimtime="00:00:27.89" resultid="5548" heatid="4800" lane="2" />
                <RESULT eventid="4425" points="484" swimtime="00:00:27.70" resultid="5554" heatid="4808" lane="2" />
                <RESULT eventid="4429" points="353" swimtime="00:00:31.28" resultid="5590" heatid="4860" lane="6" />
                <RESULT eventid="10332" points="465" swimtime="00:00:26.02" resultid="10362" heatid="10360" lane="8" entrytime="00:00:26.17" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Barbara" lastname="Campagnoli" birthdate="2009-04-13" gender="F" nation="BRA" license="366915" swrid="5600128" athleteid="1349" externalid="366915" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="494" swimtime="00:00:30.84" resultid="1350" heatid="4662" lane="1" />
                <RESULT eventid="1077" points="483" swimtime="00:00:32.18" resultid="1351" heatid="4722" lane="3" entrytime="00:00:31.78" entrycourse="SCM" />
                <RESULT eventid="1165" points="514" swimtime="00:01:08.51" resultid="1352" heatid="4914" lane="3" entrytime="00:01:13.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="475" swimtime="00:01:04.39" resultid="1353" heatid="4933" lane="2" entrytime="00:01:02.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="481" swimtime="00:00:29.25" resultid="1354" heatid="5097" lane="1" entrytime="00:00:29.31" entrycourse="SCM" />
                <RESULT eventid="1301" points="364" swimtime="00:00:39.71" resultid="1355" heatid="5031" lane="4" />
                <RESULT eventid="4411" points="487" swimtime="00:00:30.97" resultid="5336" heatid="4686" lane="2" />
                <RESULT eventid="4413" points="464" swimtime="00:00:31.48" resultid="5342" heatid="4694" lane="2" />
                <RESULT eventid="4417" points="443" swimtime="00:00:33.12" resultid="5446" heatid="4737" lane="2" />
                <RESULT eventid="4419" points="495" swimtime="00:00:31.91" resultid="5452" heatid="4745" lane="2" />
                <RESULT eventid="5801" points="366" swimtime="00:00:39.63" resultid="10163" heatid="6074" lane="3" />
                <RESULT eventid="5804" points="498" swimtime="00:00:28.92" resultid="10213" heatid="6060" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Campagnoli" birthdate="2013-03-13" gender="M" nation="BRA" license="370651" swrid="5602519" athleteid="1377" externalid="370651" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="275" swimtime="00:00:33.41" resultid="1378" heatid="4778" lane="5" entrytime="00:00:34.80" entrycourse="SCM" />
                <RESULT eventid="1105" points="227" swimtime="00:00:36.22" resultid="1379" heatid="4839" lane="2" entrytime="00:00:35.86" entrycourse="SCM" />
                <RESULT eventid="1237" points="227" swimtime="00:01:18.27" resultid="1380" heatid="4972" lane="3" entrytime="00:01:20.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="273" swimtime="00:01:09.04" resultid="1381" heatid="5006" lane="4" entrytime="00:01:12.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="219" swimtime="00:00:41.39" resultid="1383" heatid="5139" lane="3" />
                <RESULT eventid="4423" points="205" swimtime="00:00:36.87" resultid="5481" heatid="4792" lane="1" />
                <RESULT eventid="4429" points="192" swimtime="00:00:38.28" resultid="5511" heatid="4852" lane="1" />
                <RESULT eventid="5807" points="221" swimtime="00:00:41.26" resultid="10270" heatid="6036" lane="5" />
                <RESULT eventid="10332" points="284" swimtime="00:00:30.65" resultid="10363" heatid="10355" lane="1" entrytime="00:00:31.16" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Delinski" birthdate="2009-11-28" gender="F" nation="BRA" license="385190" swrid="5600150" athleteid="1356" externalid="385190" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="334" swimtime="00:00:35.12" resultid="1357" heatid="4659" lane="3" />
                <RESULT eventid="1077" points="283" swimtime="00:00:38.44" resultid="1358" heatid="4710" lane="1" />
                <RESULT eventid="1129" points="374" swimtime="00:01:26.53" resultid="1359" heatid="4887" lane="6" entrytime="00:01:24.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="325" swimtime="00:03:15.71" resultid="1360" heatid="4922" lane="4" entrytime="00:03:14.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.75" />
                    <SPLIT distance="100" swimtime="00:01:35.23" />
                    <SPLIT distance="150" swimtime="00:02:26.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="327" swimtime="00:00:33.25" resultid="1361" heatid="5085" lane="5" />
                <RESULT eventid="1301" points="400" swimtime="00:00:38.48" resultid="1362" heatid="5044" lane="3" entrytime="00:00:38.70" entrycourse="SCM" />
                <RESULT eventid="5801" points="384" swimtime="00:00:39.00" resultid="10162" heatid="6074" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Pontes Mattioli" birthdate="2011-09-10" gender="F" nation="BRA" license="366914" swrid="5602572" athleteid="1384" externalid="366914" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="320" swimtime="00:00:35.62" resultid="1385" heatid="4669" lane="6" entrytime="00:00:39.15" entrycourse="SCM" />
                <RESULT eventid="1077" points="345" swimtime="00:00:36.00" resultid="1386" heatid="4720" lane="5" entrytime="00:00:37.97" entrycourse="SCM" />
                <RESULT eventid="1165" points="339" swimtime="00:01:18.66" resultid="1387" heatid="4913" lane="5" entrytime="00:01:24.89" entrycourse="SCM" />
                <RESULT eventid="1189" points="380" swimtime="00:01:09.33" resultid="1388" heatid="4925" lane="2" />
                <RESULT eventid="1314" points="350" swimtime="00:00:32.52" resultid="1389" heatid="5090" lane="8" entrytime="00:00:33.22" entrycourse="SCM" />
                <RESULT eventid="1301" points="248" swimtime="00:00:45.15" resultid="1390" heatid="5033" lane="2" />
                <RESULT eventid="4411" points="323" swimtime="00:00:35.50" resultid="5357" heatid="4682" lane="5" />
                <RESULT eventid="4417" points="362" swimtime="00:00:35.41" resultid="5428" heatid="4733" lane="3" />
                <RESULT eventid="4419" points="311" swimtime="00:00:37.24" resultid="5435" heatid="4743" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="APAN/PONTA GROSSA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1087" status="WDR" swimtime="00:00:00.00" resultid="1402" heatid="4747" lane="3" />
                <RESULT eventid="1324" status="DNS" swimtime="00:00:00.00" resultid="5250" heatid="5122" lane="4" />
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="13038" nation="BRA" region="PR" clubid="1805" swrid="93759" name="Associação De Pais E Atletas De Natação Ws/Crb" shortname="Apan/Ws">
          <ATHLETES>
            <ATHLETE firstname="Henrique" lastname="Ueda Pritzsche" birthdate="2012-02-07" gender="M" nation="BRA" license="417110" swrid="5756912" athleteid="1917" externalid="417110" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="227" swimtime="00:00:35.61" resultid="1918" heatid="4766" lane="1" />
                <RESULT eventid="1105" points="187" swimtime="00:00:38.60" resultid="1919" heatid="4828" lane="1" />
                <RESULT eventid="1249" points="186" swimtime="00:01:24.54" resultid="1920" heatid="4980" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="220" swimtime="00:01:14.20" resultid="1921" heatid="5000" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="115" swimtime="00:00:51.25" resultid="1923" heatid="5144" lane="3" />
                <RESULT eventid="10332" points="257" swimtime="00:00:31.68" resultid="10383" heatid="10346" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Bernardi Iurk" birthdate="2012-04-14" gender="M" nation="BRA" license="408687" swrid="5725984" athleteid="1832" externalid="408687" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="163" swimtime="00:00:39.81" resultid="1833" heatid="4771" lane="1" />
                <RESULT eventid="1105" points="167" swimtime="00:00:40.11" resultid="1834" heatid="4835" lane="1" entrytime="00:00:46.55" entrycourse="SCM" />
                <RESULT eventid="1213" points="153" swimtime="00:01:43.16" resultid="1835" heatid="4951" lane="3" entrytime="00:01:57.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="158" swimtime="00:01:29.34" resultid="1836" heatid="4983" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10332" status="DNS" swimtime="00:00:00.00" resultid="10377" heatid="10351" lane="8" entrytime="00:00:36.08" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Dos Santos" birthdate="2013-06-26" gender="F" nation="BRA" license="387512" swrid="5588662" athleteid="1850" externalid="387512" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="183" swimtime="00:00:42.88" resultid="1851" heatid="4658" lane="1" />
                <RESULT eventid="1077" points="208" swimtime="00:00:42.56" resultid="1852" heatid="4716" lane="5" entrytime="00:00:43.99" entrycourse="SCM" />
                <RESULT eventid="1143" points="258" swimtime="00:02:53.10" resultid="1853" heatid="4894" lane="3" entrytime="00:03:04.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                    <SPLIT distance="100" swimtime="00:01:19.81" />
                    <SPLIT distance="150" swimtime="00:02:06.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="280" swimtime="00:01:16.80" resultid="1854" heatid="4928" lane="1" entrytime="00:01:26.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="299" swimtime="00:00:34.27" resultid="1855" heatid="5088" lane="3" entrytime="00:00:35.76" entrycourse="SCM" />
                <RESULT eventid="1301" points="88" swimtime="00:01:03.61" resultid="1856" heatid="5031" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Cravcenco Marcondes" birthdate="2011-05-06" gender="M" nation="BRA" license="406867" swrid="5723023" athleteid="1884" externalid="406867" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="272" swimtime="00:00:33.54" resultid="1885" heatid="4777" lane="3" entrytime="00:00:36.16" entrycourse="SCM" />
                <RESULT eventid="1105" points="200" swimtime="00:00:37.80" resultid="1886" heatid="4825" lane="5" />
                <RESULT eventid="1249" points="190" swimtime="00:01:23.94" resultid="1887" heatid="4982" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="278" swimtime="00:01:08.65" resultid="1888" heatid="5000" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="158" swimtime="00:00:46.11" resultid="1890" heatid="5146" lane="5" />
                <RESULT eventid="10332" points="292" swimtime="00:00:30.38" resultid="10381" heatid="10355" lane="6" entrytime="00:00:31.46" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Cravcenco Marcondes" birthdate="2012-06-23" gender="F" nation="BRA" license="406866" swrid="5725987" athleteid="1877" externalid="406866" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="139" swimtime="00:00:47.05" resultid="1878" heatid="4664" lane="3" />
                <RESULT eventid="1077" points="210" swimtime="00:00:42.45" resultid="1879" heatid="4716" lane="1" entrytime="00:00:44.16" entrycourse="SCM" />
                <RESULT eventid="1129" points="205" swimtime="00:01:45.76" resultid="1880" heatid="4885" lane="6" entrytime="00:01:53.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="193" swimtime="00:03:52.85" resultid="1881" heatid="4921" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.55" />
                    <SPLIT distance="100" swimtime="00:01:52.44" />
                    <SPLIT distance="150" swimtime="00:02:54.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="237" swimtime="00:00:37.04" resultid="1882" heatid="5085" lane="1" />
                <RESULT eventid="1301" points="196" swimtime="00:00:48.83" resultid="1883" heatid="5041" lane="6" entrytime="00:00:48.19" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Iasmim" lastname="Ferenczuk" birthdate="2013-06-06" gender="F" nation="BRA" license="414654" swrid="5755335" athleteid="1905" externalid="414654" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" status="DNS" swimtime="00:00:00.00" resultid="1906" heatid="4659" lane="2" />
                <RESULT eventid="1077" points="122" swimtime="00:00:50.78" resultid="1907" heatid="4713" lane="3" />
                <RESULT eventid="1314" points="146" swimtime="00:00:43.46" resultid="1908" heatid="5084" lane="7" />
                <RESULT eventid="1301" points="161" swimtime="00:00:52.10" resultid="1909" heatid="5032" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Daniele Silva" birthdate="2010-07-06" gender="F" nation="BRA" license="359593" swrid="5588628" athleteid="1813" externalid="359593" level="CLBO">
              <RESULTS>
                <RESULT eventid="1119" points="385" swimtime="00:02:43.38" resultid="1814" heatid="4876" lane="3" entrytime="00:02:39.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.20" />
                    <SPLIT distance="100" swimtime="00:01:19.14" />
                    <SPLIT distance="150" swimtime="00:02:01.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="379" swimtime="00:01:15.84" resultid="1815" heatid="4914" lane="4" entrytime="00:01:15.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="463" swimtime="00:01:04.91" resultid="1816" heatid="4933" lane="5" entrytime="00:01:03.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="470" swimtime="00:00:29.48" resultid="1817" heatid="5097" lane="5" entrytime="00:00:29.01" entrycourse="SCM" />
                <RESULT eventid="1301" points="363" swimtime="00:00:39.74" resultid="1818" heatid="5045" lane="7" entrytime="00:00:42.08" entrycourse="SCM" />
                <RESULT eventid="5801" points="365" swimtime="00:00:39.67" resultid="10106" heatid="6072" lane="4" />
                <RESULT eventid="5804" points="463" swimtime="00:00:29.62" resultid="10206" heatid="6058" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Reis" birthdate="2008-04-07" gender="F" nation="BRA" license="378820" swrid="5600243" athleteid="1838" externalid="378820" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="219" swimtime="00:00:40.43" resultid="1839" heatid="4667" lane="5" entrytime="00:00:44.10" entrycourse="SCM" />
                <RESULT eventid="1077" points="224" swimtime="00:00:41.55" resultid="1840" heatid="4716" lane="2" entrytime="00:00:43.66" entrycourse="SCM" />
                <RESULT eventid="1165" points="233" swimtime="00:01:29.16" resultid="1841" heatid="4906" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="267" swimtime="00:01:17.99" resultid="1842" heatid="4928" lane="4" entrytime="00:01:22.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" status="DNS" swimtime="00:00:00.00" resultid="1843" heatid="5088" lane="7" entrytime="00:00:36.88" entrycourse="SCM" />
                <RESULT eventid="1301" status="DNS" swimtime="00:00:00.00" resultid="1844" heatid="5033" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Da Reginalda" birthdate="2012-11-09" gender="M" nation="BRA" license="400275" swrid="5717253" athleteid="1864" externalid="400275" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="248" swimtime="00:00:34.60" resultid="1865" heatid="4775" lane="2" entrytime="00:00:41.92" entrycourse="SCM" />
                <RESULT eventid="1105" points="206" swimtime="00:00:37.38" resultid="1866" heatid="4838" lane="1" entrytime="00:00:37.59" entrycourse="SCM" />
                <RESULT eventid="1249" points="249" swimtime="00:01:16.72" resultid="1867" heatid="4984" lane="4" entrytime="00:01:33.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="286" swimtime="00:01:08.03" resultid="1868" heatid="5005" lane="3" entrytime="00:01:14.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="224" swimtime="00:00:41.06" resultid="1870" heatid="5151" lane="6" entrytime="00:00:45.45" entrycourse="SCM" />
                <RESULT eventid="4423" points="233" swimtime="00:00:35.32" resultid="5495" heatid="4794" lane="3" />
                <RESULT eventid="5807" points="237" swimtime="00:00:40.28" resultid="10273" heatid="6038" lane="2" />
                <RESULT eventid="10332" points="273" swimtime="00:00:31.06" resultid="10379" heatid="10354" lane="7" entrytime="00:00:32.43" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Leopoldo Goncalves" birthdate="2015-01-10" gender="M" nation="BRA" license="417109" swrid="5756907" athleteid="1910" externalid="417109" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="93" swimtime="00:00:47.96" resultid="1911" heatid="4751" lane="6" />
                <RESULT eventid="1102" points="128" swimtime="00:00:43.83" resultid="1912" heatid="4810" lane="3" />
                <RESULT eventid="1249" points="142" swimtime="00:01:32.46" resultid="1913" heatid="4978" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="168" swimtime="00:01:21.25" resultid="1914" heatid="4998" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="85" swimtime="00:00:56.68" resultid="1916" heatid="5127" lane="7" />
                <RESULT eventid="4421" points="97" swimtime="00:00:47.20" resultid="5468" heatid="4760" lane="6" />
                <RESULT eventid="4427" points="145" swimtime="00:00:42.04" resultid="5501" heatid="4821" lane="3" />
                <RESULT eventid="10329" points="187" swimtime="00:00:35.23" resultid="10382" heatid="10341" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="De Reginalda" birthdate="2011-07-22" gender="M" nation="BRA" license="400323" swrid="5717257" athleteid="1857" externalid="400323" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="350" swimtime="00:00:30.85" resultid="1858" heatid="4773" lane="4" />
                <RESULT eventid="1105" points="330" swimtime="00:00:31.97" resultid="1859" heatid="4841" lane="6" entrytime="00:00:31.54" entrycourse="SCM" />
                <RESULT eventid="1249" points="316" swimtime="00:01:10.89" resultid="1860" heatid="4986" lane="5" entrytime="00:01:09.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="406" swimtime="00:01:00.53" resultid="1861" heatid="5008" lane="6" entrytime="00:01:06.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="181" swimtime="00:00:44.09" resultid="1863" heatid="5143" lane="1" />
                <RESULT eventid="4423" points="360" swimtime="00:00:30.56" resultid="5532" heatid="4796" lane="4" />
                <RESULT eventid="4429" points="334" swimtime="00:00:31.85" resultid="5567" heatid="4856" lane="2" />
                <RESULT eventid="4431" points="251" swimtime="00:00:35.05" resultid="5573" heatid="4866" lane="2" />
                <RESULT eventid="10332" points="438" swimtime="00:00:26.53" resultid="10378" heatid="10358" lane="3" entrytime="00:00:27.61" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Bernardi Iurk" birthdate="2012-04-14" gender="M" nation="BRA" license="406940" swrid="5717245" athleteid="1826" externalid="406940" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="186" swimtime="00:00:38.10" resultid="1827" heatid="4770" lane="6" />
                <RESULT eventid="1105" points="131" swimtime="00:00:43.43" resultid="1828" heatid="4835" lane="2" entrytime="00:00:44.79" entrycourse="SCM" />
                <RESULT eventid="1227" points="242" swimtime="00:02:39.27" resultid="1829" heatid="4966" lane="6" entrytime="00:03:34.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                    <SPLIT distance="100" swimtime="00:01:17.65" />
                    <SPLIT distance="150" swimtime="00:02:00.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="252" swimtime="00:01:10.95" resultid="1830" heatid="5004" lane="4" entrytime="00:01:19.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10332" status="DNS" swimtime="00:00:00.00" resultid="10376" heatid="10352" lane="1" entrytime="00:00:34.65" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabelly" lastname="Mendonca Bello" birthdate="2008-04-15" gender="F" nation="BRA" license="376996" swrid="5600217" athleteid="1819" externalid="376996" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="363" swimtime="00:00:34.15" resultid="1820" heatid="4659" lane="6" />
                <RESULT eventid="1077" points="344" swimtime="00:00:36.03" resultid="1821" heatid="4709" lane="3" />
                <RESULT comment="SW 7.1 - Mais de uma pernada de borboleta antes da primeira pernada de peito após o início ou a virada., Na volta dos 25m." eventid="1129" status="DSQ" swimtime="00:01:23.42" resultid="1822" heatid="4886" lane="3" entrytime="00:01:24.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="465" swimtime="00:01:04.86" resultid="1823" heatid="4925" lane="6" />
                <RESULT eventid="1314" points="453" swimtime="00:00:29.84" resultid="1824" heatid="5096" lane="2" entrytime="00:00:30.61" entrycourse="SCM" />
                <RESULT eventid="1301" points="400" swimtime="00:00:38.49" resultid="1825" heatid="5044" lane="4" entrytime="00:00:38.83" entrycourse="SCM" />
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente., Na volta dos 25m." eventid="4411" status="DSQ" swimtime="00:00:35.01" resultid="5346" heatid="4688" lane="3" />
                <RESULT eventid="4417" points="350" swimtime="00:00:35.82" resultid="5456" heatid="4739" lane="3" />
                <RESULT eventid="5801" points="403" swimtime="00:00:38.38" resultid="10167" heatid="6076" lane="1" />
                <RESULT eventid="5804" points="444" swimtime="00:00:30.04" resultid="10217" heatid="6062" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leon" lastname="Bernardo Bello" birthdate="2014-11-23" gender="M" nation="BRA" license="400324" swrid="5717246" athleteid="1871" externalid="400324" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" status="DNS" swimtime="00:00:00.00" resultid="1872" heatid="4750" lane="4" />
                <RESULT eventid="1102" status="DNS" swimtime="00:00:00.00" resultid="1873" heatid="4816" lane="3" entrytime="00:00:43.70" entrycourse="SCM" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="1874" heatid="5003" lane="1" entrytime="00:01:30.44" entrycourse="SCM" />
                <RESULT eventid="1326" status="DNS" swimtime="00:00:00.00" resultid="1876" heatid="5128" lane="8" entrytime="00:00:56.63" entrycourse="SCM" />
                <RESULT eventid="10329" status="DNS" swimtime="00:00:00.00" resultid="10380" heatid="10343" lane="7" entrytime="00:00:39.54" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marjori" lastname="Leticia Oliveira" birthdate="2011-05-23" gender="F" nation="BRA" license="406869" swrid="5717279" athleteid="1898" externalid="406869" level="CLBO">
              <RESULTS>
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente., Na chegada." eventid="1064" status="DSQ" swimtime="00:00:42.65" resultid="1899" heatid="4662" lane="5" />
                <RESULT eventid="1077" points="223" swimtime="00:00:41.62" resultid="1900" heatid="4717" lane="6" entrytime="00:00:42.41" entrycourse="SCM" />
                <RESULT comment="SW 6.4 - Não tocou a borda durante a virada., Na volta dos 75m." eventid="1165" status="DSQ" swimtime="00:01:29.72" resultid="1901" heatid="4909" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="248" swimtime="00:01:19.88" resultid="1902" heatid="4925" lane="5" />
                <RESULT eventid="1314" points="288" swimtime="00:00:34.71" resultid="1903" heatid="5089" lane="5" entrytime="00:00:35.24" entrycourse="SCM" />
                <RESULT eventid="1301" points="141" swimtime="00:00:54.43" resultid="1904" heatid="5034" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cecilia" lastname="Gramms Dallarosa" birthdate="2015-01-14" gender="F" nation="BRA" license="406868" swrid="5717270" athleteid="1891" externalid="406868" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="61" swimtime="00:01:01.88" resultid="1892" heatid="4645" lane="3" />
                <RESULT eventid="1074" points="93" swimtime="00:00:55.69" resultid="1893" heatid="4699" lane="6" entrytime="00:00:56.92" entrycourse="SCM" />
                <RESULT eventid="1165" points="100" swimtime="00:01:58.07" resultid="1894" heatid="4906" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="98" swimtime="00:01:48.78" resultid="1895" heatid="4926" lane="3" entrytime="00:01:46.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="87" swimtime="00:01:03.86" resultid="1896" heatid="5021" lane="4" entrytime="00:01:06.34" entrycourse="SCM" />
                <RESULT eventid="1311" points="140" swimtime="00:00:44.14" resultid="1897" heatid="5073" lane="2" entrytime="00:00:44.22" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonia" lastname="Adam  Fracaro" birthdate="2010-04-27" gender="F" nation="BRA" license="382212" swrid="5588512" athleteid="1806" externalid="382212" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="214" swimtime="00:00:40.72" resultid="1807" heatid="4666" lane="1" />
                <RESULT eventid="1077" points="254" swimtime="00:00:39.82" resultid="1808" heatid="4719" lane="1" entrytime="00:00:39.53" entrycourse="SCM" />
                <RESULT eventid="1143" points="371" swimtime="00:02:33.49" resultid="1809" heatid="4895" lane="5" entrytime="00:02:35.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                    <SPLIT distance="100" swimtime="00:01:13.94" />
                    <SPLIT distance="150" swimtime="00:01:53.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="335" swimtime="00:01:12.29" resultid="1810" heatid="4931" lane="6" entrytime="00:01:12.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="330" swimtime="00:00:33.17" resultid="1811" heatid="5092" lane="7" entrytime="00:00:33.28" entrycourse="SCM" />
                <RESULT eventid="1301" points="207" swimtime="00:00:47.92" resultid="1812" heatid="5034" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Ferreira" birthdate="2012-12-29" gender="F" nation="BRA" license="382235" swrid="5602538" athleteid="1845" externalid="382235" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="299" swimtime="00:00:36.43" resultid="1846" heatid="4667" lane="4" entrytime="00:00:40.72" entrycourse="SCM" />
                <RESULT eventid="1077" points="270" swimtime="00:00:39.05" resultid="1847" heatid="4717" lane="3" entrytime="00:00:41.58" entrycourse="SCM" />
                <RESULT eventid="1314" points="337" swimtime="00:00:32.93" resultid="1848" heatid="5088" lane="1" entrytime="00:00:36.57" entrycourse="SCM" />
                <RESULT eventid="1301" points="191" swimtime="00:00:49.25" resultid="1849" heatid="5032" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="1202" nation="BRA" region="PR" clubid="2123" swrid="93770" name="Avulso (Paraná)" shortname="Avulso/Paraná">
          <ATHLETES>
            <ATHLETE firstname="Joao" lastname="Guilherme Ortega" birthdate="1999-08-05" gender="M" nation="BRA" license="383118" swrid="5603852" athleteid="2124" externalid="383118" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="356" status="EXH" swimtime="00:00:30.66" resultid="2125" heatid="4785" lane="6" />
                <RESULT eventid="1105" points="320" status="EXH" swimtime="00:00:32.32" resultid="2126" heatid="4850" lane="3" entrytime="00:00:30.98" entrycourse="SCM" />
                <RESULT eventid="1227" points="358" status="EXH" swimtime="00:02:19.89" resultid="2127" heatid="4968" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                    <SPLIT distance="100" swimtime="00:01:06.55" />
                    <SPLIT distance="150" swimtime="00:01:43.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="332" status="EXH" swimtime="00:01:09.75" resultid="2128" heatid="4989" lane="4" entrytime="00:01:06.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="359" status="EXH" swimtime="00:00:28.35" resultid="2129" heatid="5225" lane="5" entrytime="00:00:27.44" entrycourse="SCM" />
                <RESULT eventid="1329" points="276" status="EXH" swimtime="00:00:38.30" resultid="2130" heatid="5164" lane="5" entrytime="00:00:39.23" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="11303" nation="BRA" region="PR" clubid="2003" swrid="93760" name="Associação De Talentos Da Natação" shortname="Atn/Curitiba">
          <ATHLETES>
            <ATHLETE firstname="Isis" lastname="De Miranda" birthdate="2012-01-10" gender="F" nation="BRA" license="397278" swrid="5652886" athleteid="2076" externalid="397278" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="270" swimtime="00:00:37.70" resultid="2077" heatid="4669" lane="1" entrytime="00:00:39.13" entrycourse="SCM" />
                <RESULT eventid="1077" points="232" swimtime="00:00:41.09" resultid="2078" heatid="4708" lane="6" />
                <RESULT eventid="1165" points="259" swimtime="00:01:26.04" resultid="2079" heatid="4910" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="206" swimtime="00:01:31.50" resultid="2080" heatid="4901" lane="1" entrytime="00:01:33.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="295" swimtime="00:00:34.43" resultid="2081" heatid="5088" lane="5" entrytime="00:00:36.44" entrycourse="SCM" />
                <RESULT eventid="1301" points="155" swimtime="00:00:52.74" resultid="2082" heatid="5031" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Iglesias Prado" birthdate="2010-06-15" gender="M" nation="BRA" license="408052" swrid="5723025" athleteid="2105" externalid="408052" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="203" swimtime="00:00:36.96" resultid="2106" heatid="4777" lane="2" entrytime="00:00:36.99" entrycourse="SCM" />
                <RESULT eventid="1105" points="229" swimtime="00:00:36.13" resultid="2107" heatid="4834" lane="5" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="2108" heatid="5006" lane="6" entrytime="00:01:13.30" entrycourse="SCM" />
                <RESULT eventid="1329" points="258" swimtime="00:00:39.17" resultid="2110" heatid="5137" lane="4" />
                <RESULT eventid="10332" points="323" swimtime="00:00:29.37" resultid="10394" heatid="10354" lane="3" entrytime="00:00:31.56" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Duarte De Almeida" birthdate="2013-12-09" gender="M" nation="BRA" license="385711" swrid="5588666" athleteid="2053" externalid="385711" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="232" swimtime="00:00:35.39" resultid="2054" heatid="4778" lane="1" entrytime="00:00:35.37" entrycourse="SCM" />
                <RESULT eventid="1105" points="149" swimtime="00:00:41.68" resultid="2055" heatid="4834" lane="1" />
                <RESULT eventid="1329" points="201" swimtime="00:00:42.57" resultid="2057" heatid="5152" lane="6" entrytime="00:00:43.55" entrycourse="SCM" />
                <RESULT eventid="4425" points="224" swimtime="00:00:35.79" resultid="5476" heatid="4804" lane="2" />
                <RESULT eventid="4423" points="241" swimtime="00:00:34.91" resultid="5482" heatid="4792" lane="2" />
                <RESULT eventid="5807" points="199" swimtime="00:00:42.72" resultid="10271" heatid="6036" lane="6" />
                <RESULT eventid="10332" points="242" swimtime="00:00:32.33" resultid="10389" heatid="10354" lane="5" entrytime="00:00:31.87" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabiana" lastname="Zaleski Dallazem" birthdate="2009-05-16" gender="F" nation="BRA" license="344287" swrid="5600279" athleteid="2004" externalid="344287" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="417" swimtime="00:00:32.62" resultid="2005" heatid="4663" lane="4" />
                <RESULT eventid="1077" points="445" swimtime="00:00:33.07" resultid="2006" heatid="4722" lane="4" entrytime="00:00:31.79" entrycourse="SCM" />
                <RESULT eventid="1314" points="442" swimtime="00:00:30.08" resultid="2007" heatid="5096" lane="4" entrytime="00:00:29.92" entrycourse="SCM" />
                <RESULT eventid="1301" points="355" swimtime="00:00:40.05" resultid="2008" heatid="5038" lane="1" />
                <RESULT eventid="4411" points="336" swimtime="00:00:35.06" resultid="5339" heatid="4686" lane="5" />
                <RESULT eventid="4417" points="416" swimtime="00:00:33.80" resultid="5447" heatid="4737" lane="3" />
                <RESULT eventid="4419" points="489" swimtime="00:00:32.04" resultid="5453" heatid="4745" lane="3" />
                <RESULT eventid="5804" points="434" swimtime="00:00:30.27" resultid="10214" heatid="6060" lane="4" />
                <RESULT eventid="5801" points="349" swimtime="00:00:40.26" resultid="10327" heatid="6074" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Muller" birthdate="2009-10-10" gender="F" nation="BRA" license="376952" swrid="5600221" athleteid="2035" externalid="376952" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="331" swimtime="00:00:35.22" resultid="2036" heatid="4664" lane="1" />
                <RESULT eventid="1077" points="266" swimtime="00:00:39.26" resultid="2037" heatid="4708" lane="1" />
                <RESULT eventid="1129" points="445" swimtime="00:01:21.65" resultid="2038" heatid="4887" lane="2" entrytime="00:01:21.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="363" swimtime="00:00:32.13" resultid="2039" heatid="5094" lane="1" entrytime="00:00:31.23" entrycourse="SCM" />
                <RESULT eventid="1301" points="423" swimtime="00:00:37.78" resultid="2040" heatid="5045" lane="2" entrytime="00:00:37.40" entrycourse="SCM" />
                <RESULT eventid="5801" points="437" swimtime="00:00:37.38" resultid="10161" heatid="6074" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Bortoleto" birthdate="2008-09-05" gender="M" nation="BRA" license="406709" swrid="5717249" athleteid="2083" externalid="406709" level="CLBO">
              <RESULTS>
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente., Na volta dos 25m." eventid="1092" status="DSQ" swimtime="00:00:29.30" resultid="2084" heatid="4779" lane="4" entrytime="00:00:31.54" entrycourse="SCM" />
                <RESULT eventid="1105" points="303" swimtime="00:00:32.89" resultid="2085" heatid="4826" lane="6" />
                <RESULT eventid="1227" points="396" swimtime="00:02:15.28" resultid="2086" heatid="4965" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.60" />
                    <SPLIT distance="100" swimtime="00:01:05.31" />
                    <SPLIT distance="150" swimtime="00:01:41.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="437" swimtime="00:00:59.06" resultid="2087" heatid="5009" lane="5" entrytime="00:01:01.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="223" swimtime="00:00:41.14" resultid="2089" heatid="5144" lane="1" />
                <RESULT eventid="4429" points="338" swimtime="00:00:31.72" resultid="5595" heatid="4862" lane="5" />
                <RESULT eventid="10332" points="413" swimtime="00:00:27.06" resultid="10392" heatid="10347" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Freitas Szucs" birthdate="2011-10-02" gender="M" nation="BRA" license="377272" swrid="5588708" athleteid="2023" externalid="377272" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="224" swimtime="00:00:35.77" resultid="2024" heatid="4776" lane="6" entrytime="00:00:40.48" entrycourse="SCM" />
                <RESULT eventid="1105" points="149" swimtime="00:00:41.65" resultid="2025" heatid="4832" lane="3" />
                <RESULT eventid="1273" points="231" swimtime="00:01:13.01" resultid="2026" heatid="5005" lane="6" entrytime="00:01:18.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente., Na volta dos 25m." eventid="1329" status="DSQ" swimtime="00:00:43.99" resultid="2028" heatid="5138" lane="6" />
                <RESULT eventid="10332" points="255" swimtime="00:00:31.79" resultid="10387" heatid="10351" lane="2" entrytime="00:00:35.33" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maximilian" lastname="Hock" birthdate="2016-11-20" gender="M" nation="DEU" license="408352" athleteid="2111" externalid="408352" level="CLBO">
              <RESULTS>
                <RESULT eventid="1201" points="79" swimtime="00:00:51.49" resultid="2112" heatid="4940" lane="3" entrytime="00:01:06.07" entrycourse="SCM" />
                <RESULT eventid="1225" points="70" swimtime="00:01:00.45" resultid="2113" heatid="4960" lane="3" entrytime="00:01:07.99" entrycourse="SCM" />
                <RESULT eventid="1261" points="94" swimtime="00:00:44.29" resultid="2114" heatid="4990" lane="3" entrytime="00:00:52.09" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcos" lastname="Demchuk" birthdate="2011-06-15" gender="M" nation="BRA" license="388540" swrid="5602530" athleteid="2058" externalid="388540" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="240" swimtime="00:00:34.97" resultid="2059" heatid="4765" lane="6" />
                <RESULT eventid="1105" points="166" swimtime="00:00:40.21" resultid="2060" heatid="4831" lane="2" />
                <RESULT eventid="1273" points="315" swimtime="00:01:05.86" resultid="2061" heatid="4998" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="229" swimtime="00:00:40.74" resultid="2063" heatid="5151" lane="2" entrytime="00:00:44.85" entrycourse="SCM" />
                <RESULT eventid="10332" points="332" swimtime="00:00:29.09" resultid="10390" heatid="10352" lane="7" entrytime="00:00:33.33" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Arthur Ribeiro" birthdate="2010-02-05" gender="M" nation="BRA" license="408025" swrid="5723020" athleteid="2099" externalid="408025" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="231" swimtime="00:00:35.44" resultid="2100" heatid="4765" lane="5" />
                <RESULT eventid="1105" points="214" swimtime="00:00:36.96" resultid="2101" heatid="4830" lane="2" />
                <RESULT eventid="1213" points="331" swimtime="00:01:19.91" resultid="2102" heatid="4948" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="336" swimtime="00:00:35.86" resultid="2104" heatid="5147" lane="7" />
                <RESULT eventid="5807" points="337" swimtime="00:00:35.83" resultid="10290" heatid="6042" lane="6" />
                <RESULT eventid="10332" points="296" swimtime="00:00:30.25" resultid="10393" heatid="10348" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Camila" lastname="Duarte De Almeida" birthdate="2009-11-26" gender="F" nation="BRA" license="378819" swrid="5600152" athleteid="2041" externalid="378819" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="410" swimtime="00:00:32.80" resultid="2042" heatid="4671" lane="5" entrytime="00:00:34.13" entrycourse="SCM" />
                <RESULT eventid="1077" points="296" swimtime="00:00:37.86" resultid="2043" heatid="4712" lane="6" />
                <RESULT eventid="1314" points="425" swimtime="00:00:30.48" resultid="2044" heatid="5097" lane="7" entrytime="00:00:30.34" entrycourse="SCM" />
                <RESULT eventid="1301" points="279" swimtime="00:00:43.41" resultid="2045" heatid="5044" lane="6" entrytime="00:00:42.60" entrycourse="SCM" />
                <RESULT eventid="4411" points="393" swimtime="00:00:33.27" resultid="5340" heatid="4686" lane="6" />
                <RESULT eventid="4417" points="363" swimtime="00:00:35.39" resultid="5449" heatid="4737" lane="5" />
                <RESULT eventid="5801" points="291" swimtime="00:00:42.80" resultid="10166" heatid="6074" lane="6" />
                <RESULT eventid="5804" points="412" swimtime="00:00:30.80" resultid="10215" heatid="6060" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Guedes Braga" birthdate="2013-04-09" gender="F" nation="BRA" license="385009" swrid="5602534" athleteid="2046" externalid="385009" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="170" swimtime="00:00:43.97" resultid="2047" heatid="4666" lane="3" entrytime="00:00:46.97" entrycourse="SCM" />
                <RESULT eventid="1077" points="223" swimtime="00:00:41.63" resultid="2048" heatid="4717" lane="1" entrytime="00:00:42.39" entrycourse="SCM" />
                <RESULT eventid="1165" points="234" swimtime="00:01:28.95" resultid="2049" heatid="4912" lane="4" entrytime="00:01:33.80" entrycourse="SCM" />
                <RESULT eventid="1189" points="255" swimtime="00:01:19.22" resultid="2050" heatid="4930" lane="5" entrytime="00:01:14.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="291" swimtime="00:00:34.60" resultid="2051" heatid="5090" lane="3" entrytime="00:00:33.55" entrycourse="SCM" />
                <RESULT eventid="1301" points="136" swimtime="00:00:55.11" resultid="2052" heatid="5034" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Faria Del Valle" birthdate="2009-08-28" gender="M" nation="BRA" license="376328" swrid="5600155" athleteid="2029" externalid="376328" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="390" swimtime="00:00:29.76" resultid="2030" heatid="4774" lane="2" />
                <RESULT eventid="1105" points="329" swimtime="00:00:32.02" resultid="2031" heatid="4841" lane="1" entrytime="00:00:31.32" entrycourse="SCM" />
                <RESULT eventid="1213" status="DNS" swimtime="00:00:00.00" resultid="2032" heatid="4954" lane="1" entrytime="00:01:18.39" entrycourse="SCM" />
                <RESULT eventid="1329" points="408" swimtime="00:00:33.63" resultid="2034" heatid="5155" lane="2" entrytime="00:00:33.04" entrycourse="SCM" />
                <RESULT eventid="4423" points="358" swimtime="00:00:30.62" resultid="5552" heatid="4800" lane="6" />
                <RESULT eventid="5807" points="419" swimtime="00:00:33.34" resultid="10298" heatid="6044" lane="7" />
                <RESULT eventid="10332" points="475" swimtime="00:00:25.82" resultid="10388" heatid="10360" lane="5" entrytime="00:00:25.18" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Castellano Purkot" birthdate="2010-01-25" gender="M" nation="BRA" license="392484" swrid="5622268" athleteid="2071" externalid="392484" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="185" swimtime="00:00:38.11" resultid="2072" heatid="4768" lane="2" />
                <RESULT eventid="1105" points="221" swimtime="00:00:36.55" resultid="2073" heatid="4838" lane="3" entrytime="00:00:36.79" entrycourse="SCM" />
                <RESULT eventid="1329" points="239" swimtime="00:00:40.20" resultid="2075" heatid="5142" lane="6" />
                <RESULT eventid="10332" points="290" swimtime="00:00:30.45" resultid="10391" heatid="10356" lane="6" entrytime="00:00:29.84" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Zaleski Dallazem" birthdate="2009-05-16" gender="M" nation="BRA" license="344286" swrid="5600280" athleteid="2016" externalid="344286" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="420" swimtime="00:00:29.03" resultid="2017" heatid="4764" lane="4" />
                <RESULT eventid="1105" points="310" swimtime="00:00:32.66" resultid="2018" heatid="4828" lane="6" />
                <RESULT eventid="1213" points="404" swimtime="00:01:14.77" resultid="2019" heatid="4954" lane="4" entrytime="00:01:15.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="425" swimtime="00:00:59.61" resultid="2020" heatid="5009" lane="3" entrytime="00:01:00.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="386" swimtime="00:00:34.24" resultid="2022" heatid="5155" lane="1" entrytime="00:00:34.28" entrycourse="SCM" />
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida." eventid="4423" status="DSQ" swimtime="00:00:28.77" resultid="5551" heatid="4800" lane="5" />
                <RESULT eventid="10332" points="403" swimtime="00:00:27.29" resultid="10386" heatid="10358" lane="5" entrytime="00:00:27.90" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Manuela Souza" birthdate="2016-07-07" gender="F" nation="BRA" license="406759" swrid="5717282" athleteid="2090" externalid="406759" level="CLBO">
              <RESULTS>
                <RESULT eventid="1117" points="78" swimtime="00:00:59.07" resultid="2091" heatid="4872" lane="3" entrytime="00:01:08.54" entrycourse="SCM" />
                <RESULT eventid="1141" points="109" swimtime="00:00:59.23" resultid="2092" heatid="4891" lane="3" entrytime="00:01:10.38" entrycourse="SCM" />
                <RESULT eventid="1177" points="78" swimtime="00:00:53.64" resultid="2093" heatid="4918" lane="3" entrytime="00:01:05.10" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Kerppers Kreia" birthdate="2006-12-01" gender="M" nation="BRA" license="366815" swrid="5600195" athleteid="2009" externalid="366815" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="413" swimtime="00:00:29.19" resultid="2010" heatid="4780" lane="1" entrytime="00:00:30.33" entrycourse="SCM" />
                <RESULT eventid="1105" points="277" swimtime="00:00:33.90" resultid="2011" heatid="4826" lane="1" />
                <RESULT eventid="1227" points="513" swimtime="00:02:04.11" resultid="2012" heatid="4967" lane="2" entrytime="00:02:07.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.36" />
                    <SPLIT distance="100" swimtime="00:00:58.82" />
                    <SPLIT distance="150" swimtime="00:01:30.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="500" swimtime="00:00:56.46" resultid="2013" heatid="5011" lane="6" entrytime="00:00:57.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="258" swimtime="00:00:39.17" resultid="2015" heatid="5142" lane="7" />
                <RESULT eventid="10332" points="434" swimtime="00:00:26.62" resultid="10385" heatid="10359" lane="5" entrytime="00:00:26.26" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Neves Vianna" birthdate="2007-12-30" gender="F" nation="BRA" license="391106" swrid="5600223" athleteid="2064" externalid="391106" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="162" swimtime="00:00:44.68" resultid="2065" heatid="4659" lane="4" />
                <RESULT eventid="1077" points="203" swimtime="00:00:42.92" resultid="2066" heatid="4716" lane="4" entrytime="00:00:43.38" entrycourse="SCM" />
                <RESULT eventid="1165" points="223" swimtime="00:01:30.50" resultid="2067" heatid="4912" lane="3" entrytime="00:01:29.43" entrycourse="SCM" />
                <RESULT eventid="1189" points="234" swimtime="00:01:21.48" resultid="2068" heatid="4930" lane="6" entrytime="00:01:17.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="254" swimtime="00:00:36.16" resultid="2069" heatid="5088" lane="4" entrytime="00:00:35.96" entrycourse="SCM" />
                <RESULT eventid="1301" points="121" swimtime="00:00:57.31" resultid="2070" heatid="5038" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Goncalves Ghion" birthdate="2014-10-15" gender="F" nation="BRA" license="406912" swrid="5717269" athleteid="2094" externalid="406912" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="116" swimtime="00:00:49.92" resultid="2095" heatid="4646" lane="4" />
                <RESULT eventid="1074" points="119" swimtime="00:00:51.28" resultid="2096" heatid="4699" lane="1" entrytime="00:00:55.30" entrycourse="SCM" />
                <RESULT eventid="1298" points="139" swimtime="00:00:54.73" resultid="2097" heatid="5023" lane="5" entrytime="00:00:58.86" entrycourse="SCM" />
                <RESULT eventid="1311" points="159" swimtime="00:00:42.31" resultid="2098" heatid="5073" lane="3" entrytime="00:00:42.90" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="ATN/CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1115" points="316" status="EXH" swimtime="00:04:23.18" resultid="2117" heatid="4871" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                    <SPLIT distance="100" swimtime="00:00:59.39" />
                    <SPLIT distance="150" swimtime="00:01:35.15" />
                    <SPLIT distance="200" swimtime="00:02:10.35" />
                    <SPLIT distance="250" swimtime="00:02:44.37" />
                    <SPLIT distance="300" swimtime="00:03:22.81" />
                    <SPLIT distance="350" swimtime="00:03:48.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2053" number="1" />
                    <RELAYPOSITION athleteid="2023" number="2" />
                    <RELAYPOSITION athleteid="2071" number="3" />
                    <RELAYPOSITION athleteid="2029" number="4" />
                    <RELAYPOSITION athleteid="2083" number="5" />
                    <RELAYPOSITION athleteid="2009" number="6" />
                    <RELAYPOSITION athleteid="2058" number="7" />
                    <RELAYPOSITION athleteid="2099" number="8" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1339" points="369" status="EXH" swimtime="00:03:47.96" resultid="2118" heatid="5246" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.98" />
                    <SPLIT distance="100" swimtime="00:00:56.79" />
                    <SPLIT distance="150" swimtime="00:01:25.97" />
                    <SPLIT distance="200" swimtime="00:01:58.67" />
                    <SPLIT distance="250" swimtime="00:02:25.03" />
                    <SPLIT distance="300" swimtime="00:02:55.41" />
                    <SPLIT distance="350" swimtime="00:03:21.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2099" number="1" />
                    <RELAYPOSITION athleteid="2083" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2058" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="2053" number="4" reactiontime="0" />
                    <RELAYPOSITION athleteid="2016" number="5" reactiontime="0" />
                    <RELAYPOSITION athleteid="2071" number="6" reactiontime="0" />
                    <RELAYPOSITION athleteid="2029" number="7" reactiontime="0" />
                    <RELAYPOSITION athleteid="2009" number="8" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="ATN/CURITIBA &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1115" status="WDR" swimtime="00:00:00.00" resultid="2121" heatid="4870" lane="3" />
                <RESULT eventid="1339" status="WDR" swimtime="00:00:00.00" resultid="2122" heatid="5246" lane="7">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="2" reactiontime="0" />
                    <RELAYPOSITION number="3" reactiontime="0" />
                    <RELAYPOSITION number="4" reactiontime="0" />
                    <RELAYPOSITION number="5" reactiontime="0" />
                    <RELAYPOSITION number="6" reactiontime="0" />
                    <RELAYPOSITION number="7" reactiontime="0" />
                    <RELAYPOSITION number="8" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="ATN/CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1087" status="WDR" swimtime="00:00:00.00" resultid="2115" heatid="4748" lane="6" />
                <RESULT eventid="1324" status="DNS" swimtime="00:00:00.00" resultid="2116" heatid="5122" lane="3" />
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="ATN/CURITIBA &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1087" status="WDR" swimtime="00:00:00.00" resultid="2119" heatid="4748" lane="1" />
                <RESULT comment="SW 10.12 - Os pés perderam contato com a plataforma de partida antes que o colega de equipe anterior tocasse a borda." eventid="1324" status="DSQ" swimtime="00:04:47.97" resultid="2120" heatid="5123" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                    <SPLIT distance="100" swimtime="00:01:13.39" />
                    <SPLIT distance="150" swimtime="00:01:46.45" />
                    <SPLIT distance="200" swimtime="00:02:15.68" />
                    <SPLIT distance="250" swimtime="00:03:07.47" />
                    <SPLIT distance="300" swimtime="00:03:42.17" />
                    <SPLIT distance="350" swimtime="00:04:17.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2035" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="2094" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="2076" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="2004" number="4" status="DSQ" />
                    <RELAYPOSITION athleteid="2090" number="5" status="DSQ" />
                    <RELAYPOSITION athleteid="2046" number="6" status="DSQ" />
                    <RELAYPOSITION athleteid="2064" number="7" status="DSQ" />
                    <RELAYPOSITION athleteid="2041" number="8" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="16053" nation="BRA" region="PR" clubid="3091" swrid="93777" name="Fábrica De Nadadores" shortname="Fábrica">
          <ATHLETES>
            <ATHLETE firstname="Lucas" lastname="Silveira De Almeida" birthdate="2008-07-08" gender="M" nation="BRA" license="368152" swrid="5603912" athleteid="3197" externalid="368152" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="430" swimtime="00:00:28.80" resultid="3198" heatid="4791" lane="1" entrytime="00:00:27.94" entrycourse="SCM" />
                <RESULT eventid="1105" points="298" swimtime="00:00:33.10" resultid="3199" heatid="4844" lane="6" />
                <RESULT eventid="1237" points="376" swimtime="00:01:06.19" resultid="3200" heatid="4977" lane="2" entrytime="00:01:01.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="372" swimtime="00:02:46.93" resultid="3201" heatid="4994" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                    <SPLIT distance="100" swimtime="00:01:19.27" />
                    <SPLIT distance="150" swimtime="00:02:03.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="392" swimtime="00:00:27.53" resultid="3202" heatid="5217" lane="4" />
                <RESULT eventid="1329" points="370" swimtime="00:00:34.75" resultid="3203" heatid="5157" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Garcia Saqueto" birthdate="2015-08-16" gender="M" nation="BRA" license="418300" athleteid="3480" externalid="418300" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="46" swimtime="00:01:00.40" resultid="3481" heatid="4750" lane="3" />
                <RESULT eventid="1102" points="82" swimtime="00:00:50.84" resultid="3482" heatid="4812" lane="1" />
                <RESULT eventid="1326" points="74" swimtime="00:00:59.29" resultid="3484" heatid="5126" lane="8" />
                <RESULT eventid="4427" points="81" swimtime="00:00:50.90" resultid="5504" heatid="4821" lane="5" />
                <RESULT eventid="10329" points="100" swimtime="00:00:43.40" resultid="10482" heatid="10340" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabel" lastname="Rezende" birthdate="2013-12-13" gender="F" nation="BRA" license="370657" swrid="5603900" athleteid="3127" externalid="370657" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="180" swimtime="00:00:43.16" resultid="3128" heatid="4672" lane="5" />
                <RESULT comment="SW 6.4 - Não começou a executar a virada imediatamente após virar para a posição de peito.  (Horário: 10:21)" eventid="1077" status="DSQ" swimtime="00:00:44.64" resultid="3129" heatid="4726" lane="6" entrytime="00:00:45.88" entrycourse="SCM" />
                <RESULT eventid="1165" points="186" swimtime="00:01:35.99" resultid="3130" heatid="4916" lane="3" entrytime="00:01:38.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="211" swimtime="00:01:24.28" resultid="3131" heatid="4937" lane="2" entrytime="00:01:24.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="236" swimtime="00:00:37.10" resultid="3132" heatid="5100" lane="6" entrytime="00:00:36.79" entrycourse="SCM" />
                <RESULT eventid="1301" points="171" swimtime="00:00:51.04" resultid="3133" heatid="5049" lane="5" entrytime="00:00:53.10" entrycourse="SCM" />
                <RESULT eventid="5801" points="176" swimtime="00:00:50.57" resultid="10015" heatid="6067" lane="5" />
                <RESULT eventid="5804" points="231" swimtime="00:00:37.34" resultid="10055" heatid="6053" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Bagatim" birthdate="2014-05-27" gender="F" nation="BRA" license="378353" swrid="5236649" athleteid="3225" externalid="378353" level="MRGA">
              <RESULTS>
                <RESULT eventid="1061" points="279" swimtime="00:00:37.31" resultid="3226" heatid="4654" lane="3" entrytime="00:00:37.88" entrycourse="SCM" />
                <RESULT eventid="1074" points="182" swimtime="00:00:44.52" resultid="3227" heatid="4705" lane="4" entrytime="00:00:43.27" entrycourse="SCM" />
                <RESULT eventid="1153" points="182" swimtime="00:01:35.23" resultid="3228" heatid="4902" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="249" swimtime="00:01:19.84" resultid="3229" heatid="4937" lane="3" entrytime="00:01:21.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="201" swimtime="00:00:48.40" resultid="3230" heatid="5028" lane="3" entrytime="00:00:47.79" entrycourse="SCM" />
                <RESULT eventid="1311" points="293" swimtime="00:00:34.50" resultid="3231" heatid="5079" lane="3" entrytime="00:00:34.23" entrycourse="SCM" />
                <RESULT eventid="4415" points="179" swimtime="00:00:44.79" resultid="9012" heatid="9004" lane="5" />
                <RESULT eventid="4409" points="313" swimtime="00:00:35.89" resultid="9018" heatid="9002" lane="4" />
                <RESULT eventid="4433" points="204" swimtime="00:00:48.16" resultid="10005" heatid="6065" lane="1" />
                <RESULT eventid="4439" points="271" swimtime="00:00:35.42" resultid="10044" heatid="6051" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Voltarelli Souza" birthdate="2014-07-26" gender="M" nation="BRA" license="410202" swrid="5748710" athleteid="3430" externalid="410202" level="MRGA">
              <RESULTS>
                <RESULT eventid="1089" points="113" swimtime="00:00:44.92" resultid="3431" heatid="4759" lane="1" entrytime="00:00:49.48" entrycourse="SCM" />
                <RESULT eventid="1102" points="101" swimtime="00:00:47.41" resultid="3432" heatid="4820" lane="6" entrytime="00:00:47.32" entrycourse="SCM" />
                <RESULT eventid="1213" points="140" swimtime="00:01:46.21" resultid="3433" heatid="4956" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="119" swimtime="00:01:38.17" resultid="3434" heatid="4987" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="140" swimtime="00:00:38.80" resultid="3435" heatid="5193" lane="4" entrytime="00:00:41.72" entrycourse="SCM" />
                <RESULT eventid="1326" points="124" swimtime="00:00:49.98" resultid="3436" heatid="5134" lane="1" entrytime="00:00:51.86" entrycourse="SCM" />
                <RESULT eventid="4427" points="116" swimtime="00:00:45.25" resultid="9033" heatid="9008" lane="6" />
                <RESULT eventid="4445" points="125" swimtime="00:00:49.79" resultid="10119" heatid="6035" lane="4" />
                <RESULT eventid="4451" points="144" swimtime="00:00:38.46" resultid="10233" heatid="6019" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Kenji Yamaguchi" birthdate="2011-08-25" gender="M" nation="BRA" license="385708" swrid="5603862" athleteid="3169" externalid="385708" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="318" swimtime="00:00:31.84" resultid="3170" heatid="4789" lane="2" entrytime="00:00:33.98" entrycourse="SCM" />
                <RESULT eventid="1105" points="221" swimtime="00:00:36.53" resultid="3171" heatid="4845" lane="3" />
                <RESULT eventid="1237" points="289" swimtime="00:01:12.24" resultid="3172" heatid="4976" lane="3" entrytime="00:01:14.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="260" swimtime="00:03:08.16" resultid="3173" heatid="4994" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.08" />
                    <SPLIT distance="100" swimtime="00:01:30.46" />
                    <SPLIT distance="150" swimtime="00:02:19.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="256" swimtime="00:00:31.75" resultid="3174" heatid="5221" lane="3" entrytime="00:00:32.94" entrycourse="SCM" />
                <RESULT comment="SW 7.1 - Mais de uma pernada de borboleta antes da primeira pernada de peito após o início ou a virada.  (Horário: 10:48)" eventid="1329" status="DSQ" swimtime="00:00:39.75" resultid="3175" heatid="5160" lane="6" />
                <RESULT eventid="4423" points="313" swimtime="00:00:32.00" resultid="5707" heatid="4797" lane="3" />
                <RESULT eventid="4425" points="290" swimtime="00:00:32.85" resultid="5735" heatid="4806" lane="5" />
                <RESULT eventid="4429" points="212" swimtime="00:00:37.07" resultid="5761" heatid="4857" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robsson" lastname="Tows Oliveira" birthdate="2014-03-05" gender="M" nation="BRA" license="392107" swrid="5603922" athleteid="3341" externalid="392107" level="MRGA">
              <RESULTS>
                <RESULT eventid="1089" points="92" swimtime="00:00:48.05" resultid="3342" heatid="4757" lane="4" />
                <RESULT eventid="1102" points="92" swimtime="00:00:48.90" resultid="3343" heatid="4818" lane="2" />
                <RESULT eventid="1213" points="141" swimtime="00:01:46.06" resultid="3344" heatid="4956" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="138" swimtime="00:01:26.72" resultid="3345" heatid="5014" lane="3" entrytime="00:01:26.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="140" swimtime="00:00:38.79" resultid="3346" heatid="5194" lane="5" entrytime="00:00:38.50" entrycourse="SCM" />
                <RESULT eventid="1326" points="136" swimtime="00:00:48.40" resultid="3347" heatid="5134" lane="4" entrytime="00:00:48.60" entrycourse="SCM" />
                <RESULT eventid="4445" points="128" swimtime="00:00:49.39" resultid="10117" heatid="6035" lane="2" />
                <RESULT eventid="4451" points="148" swimtime="00:00:38.03" resultid="10232" heatid="6019" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theodoro" lastname="Marques Serra" birthdate="2009-11-24" gender="M" nation="BRA" license="370661" swrid="5603870" athleteid="3155" externalid="370661" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="337" swimtime="00:00:31.23" resultid="3156" heatid="4790" lane="4" entrytime="00:00:30.22" entrycourse="SCM" />
                <RESULT eventid="1105" points="226" swimtime="00:00:36.25" resultid="3157" heatid="4850" lane="2" entrytime="00:00:33.73" entrycourse="SCM" />
                <RESULT eventid="1227" points="439" swimtime="00:02:10.72" resultid="3158" heatid="5254" lane="3" entrytime="00:02:12.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                    <SPLIT distance="100" swimtime="00:01:02.19" />
                    <SPLIT distance="150" swimtime="00:01:36.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="322" swimtime="00:01:10.49" resultid="3159" heatid="4989" lane="5" entrytime="00:01:08.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="335" swimtime="00:00:29.01" resultid="3160" heatid="5225" lane="6" entrytime="00:00:27.79" entrycourse="SCM" />
                <RESULT eventid="1329" points="293" swimtime="00:00:37.56" resultid="3161" heatid="5158" lane="5" />
                <RESULT eventid="4423" points="351" swimtime="00:00:30.83" resultid="5720" heatid="4801" lane="5" />
                <RESULT eventid="4425" points="379" swimtime="00:00:30.04" resultid="5741" heatid="4808" lane="5" />
                <RESULT eventid="4429" points="313" swimtime="00:00:32.54" resultid="5768" heatid="4861" lane="3" />
                <RESULT eventid="4431" points="373" swimtime="00:00:30.71" resultid="5790" heatid="4868" lane="5" />
                <RESULT eventid="5807" points="292" swimtime="00:00:37.58" resultid="10146" heatid="6045" lane="4" />
                <RESULT eventid="5810" points="380" swimtime="00:00:27.81" resultid="10260" heatid="6029" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jennifer" lastname="De Abreu" birthdate="2009-11-07" gender="F" nation="BRA" license="356212" swrid="5600144" athleteid="3099" externalid="356212" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="436" swimtime="00:00:32.13" resultid="3100" heatid="4671" lane="4" entrytime="00:00:32.20" entrycourse="SCM" />
                <RESULT eventid="1077" points="327" swimtime="00:00:36.62" resultid="3101" heatid="4710" lane="3" />
                <RESULT eventid="1129" points="369" swimtime="00:01:26.88" resultid="3102" heatid="4884" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="349" swimtime="00:01:17.95" resultid="3103" heatid="4909" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="441" swimtime="00:00:30.11" resultid="3104" heatid="5097" lane="6" entrytime="00:00:29.61" entrycourse="SCM" />
                <RESULT eventid="1301" status="DNS" swimtime="00:00:00.00" resultid="3105" heatid="5033" lane="6" />
                <RESULT eventid="4411" points="407" swimtime="00:00:32.88" resultid="5337" heatid="4686" lane="3" />
                <RESULT eventid="4413" points="381" swimtime="00:00:33.62" resultid="5343" heatid="4694" lane="3" />
                <RESULT eventid="4417" points="339" swimtime="00:00:36.21" resultid="5448" heatid="4737" lane="4" />
                <RESULT eventid="5804" points="424" swimtime="00:00:30.50" resultid="10210" heatid="6060" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luana" lastname="Siqueira Lopes" birthdate="2012-04-28" gender="F" nation="BRA" license="414671" swrid="5755342" athleteid="3458" externalid="414671" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="272" swimtime="00:00:37.60" resultid="3459" heatid="4663" lane="5" />
                <RESULT eventid="1077" points="234" swimtime="00:00:40.95" resultid="3460" heatid="4711" lane="6" />
                <RESULT eventid="1189" points="322" swimtime="00:01:13.29" resultid="3461" heatid="4925" lane="1" />
                <RESULT eventid="1314" points="353" swimtime="00:00:32.43" resultid="3462" heatid="5083" lane="6" />
                <RESULT eventid="1301" points="191" swimtime="00:00:49.18" resultid="3463" heatid="5036" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Tiemi Yamaguchi" birthdate="2013-02-28" gender="F" nation="BRA" license="385707" swrid="5603920" athleteid="3246" externalid="385707" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="269" swimtime="00:00:37.75" resultid="3247" heatid="4676" lane="2" entrytime="00:00:37.38" entrycourse="SCM" />
                <RESULT eventid="1077" points="259" swimtime="00:00:39.60" resultid="3248" heatid="4726" lane="3" entrytime="00:00:41.67" entrycourse="SCM" />
                <RESULT eventid="1119" points="292" swimtime="00:02:59.21" resultid="3249" heatid="4877" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.56" />
                    <SPLIT distance="100" swimtime="00:01:29.69" />
                    <SPLIT distance="150" swimtime="00:02:14.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="254" swimtime="00:01:25.31" resultid="3250" heatid="4903" lane="2" entrytime="00:01:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="257" swimtime="00:00:36.06" resultid="3251" heatid="5100" lane="4" entrytime="00:00:35.18" entrycourse="SCM" />
                <RESULT eventid="1301" points="235" swimtime="00:00:45.92" resultid="3252" heatid="5050" lane="2" entrytime="00:00:46.26" entrycourse="SCM" />
                <RESULT eventid="4411" points="300" swimtime="00:00:36.38" resultid="5610" heatid="4679" lane="4" />
                <RESULT eventid="4413" points="302" swimtime="00:00:36.32" resultid="5635" heatid="4690" lane="6" />
                <RESULT eventid="4417" points="277" swimtime="00:00:38.73" resultid="5652" heatid="4730" lane="3" />
                <RESULT eventid="4419" points="281" swimtime="00:00:38.55" resultid="5678" heatid="4741" lane="5" />
                <RESULT eventid="5801" points="245" swimtime="00:00:45.31" resultid="10012" heatid="6067" lane="2" />
                <RESULT eventid="5804" points="251" swimtime="00:00:36.32" resultid="10054" heatid="6053" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Magalhães Rezende" birthdate="2010-05-29" gender="F" nation="BRA" license="366960" swrid="5588793" athleteid="3176" externalid="366960" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="270" swimtime="00:00:37.69" resultid="3177" heatid="4672" lane="1" />
                <RESULT eventid="1077" points="278" swimtime="00:00:38.68" resultid="3178" heatid="4724" lane="4" />
                <RESULT eventid="1165" points="290" swimtime="00:01:22.84" resultid="3179" heatid="4917" lane="2" entrytime="00:01:21.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="344" swimtime="00:02:37.29" resultid="3180" heatid="4897" lane="5" entrytime="00:02:37.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.08" />
                    <SPLIT distance="100" swimtime="00:01:14.79" />
                    <SPLIT distance="150" swimtime="00:01:56.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="297" swimtime="00:00:34.36" resultid="3181" heatid="5102" lane="3" entrytime="00:00:31.59" entrycourse="SCM" />
                <RESULT eventid="1301" points="283" swimtime="00:00:43.21" resultid="3182" heatid="5048" lane="1" />
                <RESULT eventid="4411" points="283" swimtime="00:00:37.11" resultid="5626" heatid="4685" lane="4" />
                <RESULT eventid="4417" points="291" swimtime="00:00:38.09" resultid="5669" heatid="4736" lane="4" />
                <RESULT eventid="4419" points="300" swimtime="00:00:37.70" resultid="5688" heatid="4744" lane="6" />
                <RESULT eventid="5801" points="301" swimtime="00:00:42.32" resultid="10027" heatid="6073" lane="1" />
                <RESULT eventid="5804" points="333" swimtime="00:00:33.07" resultid="10070" heatid="6059" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Pazinato" birthdate="2011-01-05" gender="M" nation="BRA" license="368149" swrid="5603889" athleteid="3190" externalid="368149" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="301" swimtime="00:00:32.43" resultid="3191" heatid="4782" lane="2" />
                <RESULT eventid="1105" points="243" swimtime="00:00:35.41" resultid="3192" heatid="4844" lane="1" />
                <RESULT eventid="1249" points="265" swimtime="00:01:15.20" resultid="3193" heatid="4989" lane="6" entrytime="00:01:15.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="313" swimtime="00:01:06.01" resultid="3194" heatid="5016" lane="3" entrytime="00:01:04.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="319" swimtime="00:00:29.50" resultid="3195" heatid="5223" lane="2" entrytime="00:00:29.52" entrycourse="SCM" />
                <RESULT eventid="1329" points="204" swimtime="00:00:42.35" resultid="3196" heatid="5159" lane="3" />
                <RESULT eventid="4423" points="300" swimtime="00:00:32.46" resultid="5709" heatid="4797" lane="4" />
                <RESULT eventid="4429" points="264" swimtime="00:00:34.45" resultid="5759" heatid="4857" lane="3" />
                <RESULT eventid="5807" points="205" swimtime="00:00:42.29" resultid="10136" heatid="6041" lane="4" />
                <RESULT eventid="5810" points="335" swimtime="00:00:29.01" resultid="10248" heatid="6025" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Traci Rodrigues" birthdate="2011-03-06" gender="M" nation="BRA" license="406927" swrid="5718893" athleteid="3120" externalid="406927" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="138" swimtime="00:00:42.03" resultid="3121" heatid="4784" lane="3" />
                <RESULT eventid="1105" points="118" swimtime="00:00:45.05" resultid="3122" heatid="4847" lane="3" entrytime="00:00:47.06" entrycourse="SCM" />
                <RESULT comment="SW 7.4 - Movimentos das pernas não simultâneos.  (Horário: 17:50), Durante a fase submersa dos 25m, 50m e 75m." eventid="1213" status="DSQ" swimtime="00:01:40.14" resultid="3123" heatid="4958" lane="6" entrytime="00:01:39.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="198" swimtime="00:01:16.90" resultid="3124" heatid="5012" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="205" swimtime="00:00:34.14" resultid="3125" heatid="5220" lane="3" entrytime="00:00:34.20" entrycourse="SCM" />
                <RESULT comment="SW 7.4 - Movimentos das pernas não simultâneos.  (Horário: 10:48)" eventid="1329" status="DSQ" swimtime="00:00:45.50" resultid="3126" heatid="5160" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Traci Rodrigues" birthdate="2014-10-27" gender="M" nation="BRA" license="406926" swrid="5726001" athleteid="3396" externalid="406926" level="MRGA">
              <RESULTS>
                <RESULT eventid="1089" points="44" swimtime="00:01:01.15" resultid="3397" heatid="4758" lane="6" entrytime="00:01:06.36" entrycourse="SCM" />
                <RESULT eventid="1102" points="71" swimtime="00:00:53.27" resultid="3398" heatid="4819" lane="6" />
                <RESULT eventid="1213" points="88" swimtime="00:02:04.25" resultid="3399" heatid="4956" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="105" swimtime="00:01:34.84" resultid="3400" heatid="5012" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="133" swimtime="00:00:39.40" resultid="3401" heatid="5193" lane="2" entrytime="00:00:42.21" entrycourse="SCM" />
                <RESULT eventid="1326" points="93" swimtime="00:00:55.03" resultid="3402" heatid="5133" lane="3" entrytime="00:00:55.69" entrycourse="SCM" />
                <RESULT eventid="4445" points="101" swimtime="00:00:53.44" resultid="10120" heatid="6035" lane="5" />
                <RESULT eventid="4451" points="117" swimtime="00:00:41.20" resultid="10234" heatid="6019" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Rossi" birthdate="2012-05-21" gender="M" nation="BRA" license="378346" swrid="5603901" athleteid="3218" externalid="378346" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="187" swimtime="00:00:38.03" resultid="3219" heatid="4788" lane="5" entrytime="00:00:37.07" entrycourse="SCM" />
                <RESULT eventid="1105" points="176" swimtime="00:00:39.38" resultid="3220" heatid="4849" lane="2" entrytime="00:00:38.49" entrycourse="SCM" />
                <RESULT eventid="1203" points="210" swimtime="00:02:57.59" resultid="3221" heatid="4944" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.73" />
                    <SPLIT distance="100" swimtime="00:01:26.82" />
                    <SPLIT distance="150" swimtime="00:02:13.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="258" swimtime="00:01:10.38" resultid="3222" heatid="5016" lane="5" entrytime="00:01:12.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="261" swimtime="00:00:31.54" resultid="3223" heatid="5221" lane="2" entrytime="00:00:33.12" entrycourse="SCM" />
                <RESULT eventid="1329" points="155" swimtime="00:00:46.36" resultid="3224" heatid="5159" lane="2" />
                <RESULT eventid="5807" points="171" swimtime="00:00:44.92" resultid="10132" heatid="6039" lane="6" />
                <RESULT eventid="5810" points="260" swimtime="00:00:31.58" resultid="10242" heatid="6023" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Covatti Anzoategui" birthdate="2013-04-13" gender="F" nation="BRA" license="420633" athleteid="3485" externalid="420633" level="MRGA">
              <RESULTS>
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 9:06), Na volta dos 25m." eventid="1064" status="DSQ" swimtime="00:01:11.55" resultid="3486" heatid="4672" lane="3" />
                <RESULT comment="SW 6.4 - Não começou a executar a virada imediatamente após virar para a posição de peito.  (Horário: 10:16), Na volta dos 25m." eventid="1077" status="DSQ" swimtime="00:00:53.76" resultid="3487" heatid="4724" lane="6" />
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 15:56), Na volta dos 25m." eventid="1129" status="DSQ" swimtime="00:02:07.18" resultid="3488" heatid="4888" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.98" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 6.4 - A virada não foi iniciada após a conclusão do movimento de braço, após sair da posição de costas.  (Horário: 16:26), Na volta dos 25m." eventid="1165" status="DSQ" swimtime="00:02:05.77" resultid="3489" heatid="4916" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="102" swimtime="00:00:48.96" resultid="3490" heatid="5098" lane="5" />
                <RESULT eventid="1301" points="110" swimtime="00:00:59.15" resultid="3491" heatid="5048" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="De Ormeno" birthdate="2014-04-02" gender="M" nation="BRA" license="408702" swrid="5740009" athleteid="3423" externalid="408702" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="145" swimtime="00:00:41.37" resultid="3424" heatid="4750" lane="2" />
                <RESULT eventid="1102" points="164" swimtime="00:00:40.39" resultid="3425" heatid="4817" lane="2" entrytime="00:00:40.25" entrycourse="SCM" />
                <RESULT eventid="1249" points="145" swimtime="00:01:31.82" resultid="3426" heatid="4982" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="170" swimtime="00:01:20.84" resultid="3427" heatid="5004" lane="5" entrytime="00:01:21.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="78" swimtime="00:00:58.26" resultid="3429" heatid="5126" lane="5" />
                <RESULT eventid="4421" points="150" swimtime="00:00:40.88" resultid="5471" heatid="4761" lane="3" />
                <RESULT eventid="4427" points="170" swimtime="00:00:39.91" resultid="5505" heatid="4822" lane="1" />
                <RESULT eventid="10329" status="DSQ" swimtime="00:00:34.75" resultid="10478" heatid="10345" lane="4" entrytime="00:00:34.65" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monique" lastname="Istake" birthdate="2012-04-03" gender="F" nation="BRA" license="372023" swrid="5603857" athleteid="3141" externalid="372023" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="396" swimtime="00:00:33.19" resultid="3142" heatid="4677" lane="1" entrytime="00:00:34.99" entrycourse="SCM" />
                <RESULT eventid="1077" points="269" swimtime="00:00:39.07" resultid="3143" heatid="4723" lane="4" />
                <RESULT eventid="1179" points="298" swimtime="00:03:21.38" resultid="3144" heatid="4923" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.54" />
                    <SPLIT distance="100" swimtime="00:01:37.23" />
                    <SPLIT distance="150" swimtime="00:02:30.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="318" swimtime="00:01:19.13" resultid="3145" heatid="4903" lane="5" entrytime="00:01:25.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="366" swimtime="00:00:32.05" resultid="3146" heatid="5101" lane="1" entrytime="00:00:34.12" entrycourse="SCM" />
                <RESULT eventid="1301" points="295" swimtime="00:00:42.61" resultid="3147" heatid="5050" lane="4" entrytime="00:00:44.84" entrycourse="SCM" />
                <RESULT eventid="4411" points="368" swimtime="00:00:34.02" resultid="5613" heatid="4681" lane="1" />
                <RESULT eventid="4413" points="388" swimtime="00:00:33.42" resultid="5637" heatid="4691" lane="5" />
                <RESULT eventid="4417" points="300" swimtime="00:00:37.70" resultid="5657" heatid="4732" lane="2" />
                <RESULT eventid="4419" points="306" swimtime="00:00:37.46" resultid="5681" heatid="4742" lane="5" />
                <RESULT eventid="5801" points="312" swimtime="00:00:41.80" resultid="10019" heatid="6069" lane="3" />
                <RESULT eventid="5804" points="375" swimtime="00:00:31.77" resultid="10057" heatid="6055" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="Jacobsen Donati" birthdate="2011-07-14" gender="M" nation="BRA" license="391851" swrid="5615735" athleteid="3162" externalid="391851" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="351" swimtime="00:00:30.83" resultid="3163" heatid="4786" lane="5" />
                <RESULT eventid="1105" points="348" swimtime="00:00:31.42" resultid="3164" heatid="4843" lane="2" />
                <RESULT eventid="1203" points="379" swimtime="00:02:25.95" resultid="3165" heatid="4945" lane="2" entrytime="00:02:33.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                    <SPLIT distance="100" swimtime="00:01:11.13" />
                    <SPLIT distance="150" swimtime="00:01:49.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1237" points="323" swimtime="00:01:09.61" resultid="3166" heatid="4975" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="347" swimtime="00:00:28.67" resultid="3167" heatid="5224" lane="3" entrytime="00:00:28.14" entrycourse="SCM" />
                <RESULT eventid="1329" points="193" swimtime="00:00:43.11" resultid="3168" heatid="5158" lane="6" />
                <RESULT eventid="4423" points="353" swimtime="00:00:30.75" resultid="5706" heatid="4797" lane="2" />
                <RESULT eventid="4425" points="359" swimtime="00:00:30.59" resultid="5734" heatid="4806" lane="4" />
                <RESULT eventid="4429" points="306" swimtime="00:00:32.78" resultid="5757" heatid="4857" lane="1" />
                <RESULT eventid="4431" points="363" swimtime="00:00:30.97" resultid="5783" heatid="4866" lane="4" />
                <RESULT eventid="5807" points="205" swimtime="00:00:42.31" resultid="10138" heatid="6041" lane="6" />
                <RESULT eventid="5810" points="400" swimtime="00:00:27.35" resultid="10247" heatid="6025" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elen" lastname="Torres Gomes" birthdate="2015-10-15" gender="F" nation="BRA" license="396850" swrid="5641777" athleteid="3295" externalid="396850" level="MRGA">
              <RESULTS>
                <RESULT eventid="1061" points="58" swimtime="00:01:02.76" resultid="3296" heatid="4653" lane="1" />
                <RESULT eventid="1074" points="89" swimtime="00:00:56.55" resultid="3297" heatid="4705" lane="1" entrytime="00:00:52.93" entrycourse="SCM" />
                <RESULT eventid="1129" points="86" swimtime="00:02:20.82" resultid="3298" heatid="4888" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="80" swimtime="00:01:56.44" resultid="3299" heatid="4935" lane="3" entrytime="00:02:13.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="75" swimtime="00:01:06.98" resultid="3300" heatid="5027" lane="1" entrytime="00:01:07.94" entrycourse="SCM" />
                <RESULT eventid="1311" points="89" swimtime="00:00:51.23" resultid="3301" heatid="5077" lane="3" entrytime="00:00:52.88" entrycourse="SCM" />
                <RESULT eventid="4415" points="91" swimtime="00:00:55.96" resultid="9009" heatid="9003" lane="4" />
                <RESULT eventid="4409" points="55" swimtime="00:01:04.08" resultid="9015" heatid="9001" lane="4" />
                <RESULT eventid="4433" points="90" swimtime="00:01:03.23" resultid="10002" heatid="5030" lane="2" />
                <RESULT eventid="4439" points="97" swimtime="00:00:49.80" resultid="10040" heatid="6049" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Taparo" birthdate="2012-04-20" gender="F" nation="BRA" license="407283" swrid="5688565" athleteid="3413" externalid="407283" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="172" swimtime="00:00:43.80" resultid="3414" heatid="4673" lane="1" />
                <RESULT eventid="1077" points="182" swimtime="00:00:44.53" resultid="3415" heatid="4726" lane="1" entrytime="00:00:45.66" entrycourse="SCM" />
                <RESULT eventid="1165" points="159" swimtime="00:01:41.22" resultid="3416" heatid="4915" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="220" swimtime="00:01:23.14" resultid="3417" heatid="4935" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="210" swimtime="00:00:38.52" resultid="3418" heatid="5099" lane="5" entrytime="00:00:37.59" entrycourse="SCM" />
                <RESULT comment="SW 7.1 - Mais de uma pernada de borboleta antes da primeira pernada de peito após o início ou a virada.  (Horário: 8:26), Após a largada." eventid="1301" status="DSQ" swimtime="00:00:55.61" resultid="3419" heatid="5046" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Braga" birthdate="2010-05-07" gender="M" nation="BRA" license="378345" swrid="5343953" athleteid="3092" externalid="378345" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="338" swimtime="00:00:31.22" resultid="3093" heatid="4783" lane="2" />
                <RESULT eventid="1105" points="207" swimtime="00:00:37.34" resultid="3094" heatid="4845" lane="6" />
                <RESULT eventid="1213" points="434" swimtime="00:01:13.01" resultid="3095" heatid="4959" lane="1" entrytime="00:01:12.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="444" swimtime="00:02:37.49" resultid="3096" heatid="4995" lane="3" entrytime="00:02:39.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                    <SPLIT distance="100" swimtime="00:01:17.22" />
                    <SPLIT distance="150" swimtime="00:01:57.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="277" swimtime="00:00:30.92" resultid="3097" heatid="5223" lane="4" entrytime="00:00:29.36" entrycourse="SCM" />
                <RESULT eventid="1329" points="409" swimtime="00:00:33.61" resultid="3098" heatid="5165" lane="1" entrytime="00:00:33.59" entrycourse="SCM" />
                <RESULT eventid="4423" points="325" swimtime="00:00:31.62" resultid="5713" heatid="4799" lane="1" />
                <RESULT eventid="4425" points="365" swimtime="00:00:30.42" resultid="5737" heatid="4807" lane="4" />
                <RESULT eventid="4429" points="193" swimtime="00:00:38.20" resultid="5764" heatid="4859" lane="2" />
                <RESULT eventid="4431" points="220" swimtime="00:00:36.61" resultid="5787" heatid="4867" lane="5" />
                <RESULT eventid="5807" points="434" swimtime="00:00:32.94" resultid="10140" heatid="6043" lane="1" />
                <RESULT eventid="5810" points="356" swimtime="00:00:28.43" resultid="10252" heatid="6027" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rodrigo" lastname="Zanatta Duda" birthdate="2011-09-12" gender="M" nation="BRA" license="406917" swrid="5717307" athleteid="3368" externalid="406917" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="160" swimtime="00:00:40.05" resultid="3369" heatid="4764" lane="2" />
                <RESULT eventid="1105" points="262" swimtime="00:00:34.54" resultid="3370" heatid="4837" lane="1" entrytime="00:00:39.35" entrycourse="SCM" />
                <RESULT eventid="1203" points="287" swimtime="00:02:39.98" resultid="3371" heatid="4942" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                    <SPLIT distance="100" swimtime="00:01:18.14" />
                    <SPLIT distance="150" swimtime="00:01:59.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="264" swimtime="00:01:15.29" resultid="3372" heatid="4985" lane="1" entrytime="00:01:25.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="176" swimtime="00:00:44.49" resultid="3374" heatid="5147" lane="5" />
                <RESULT eventid="4429" points="271" swimtime="00:00:34.14" resultid="5570" heatid="4856" lane="5" />
                <RESULT eventid="10332" points="263" swimtime="00:00:31.44" resultid="10475" heatid="10349" lane="8" entrytime="00:00:37.14" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Ribeiro Melo" birthdate="2013-02-25" gender="M" nation="BRA" license="406921" swrid="5717293" athleteid="3382" externalid="406921" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="112" swimtime="00:00:45.04" resultid="3383" heatid="4766" lane="5" />
                <RESULT eventid="1105" points="136" swimtime="00:00:42.99" resultid="3384" heatid="4836" lane="6" entrytime="00:00:43.35" entrycourse="SCM" />
                <RESULT eventid="1227" points="195" swimtime="00:02:51.11" resultid="3385" heatid="4962" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.05" />
                    <SPLIT distance="100" swimtime="00:01:24.49" />
                    <SPLIT distance="150" swimtime="00:02:08.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="138" swimtime="00:01:33.49" resultid="3386" heatid="4984" lane="5" entrytime="00:01:47.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="96" swimtime="00:00:54.45" resultid="3388" heatid="5148" lane="4" entrytime="00:00:55.53" entrycourse="SCM" />
                <RESULT eventid="10332" points="180" swimtime="00:00:35.68" resultid="10476" heatid="10350" lane="3" entrytime="00:00:35.86" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Borges Duarte" birthdate="2014-02-10" gender="F" nation="BRA" license="408688" swrid="5725985" athleteid="3420" externalid="408688" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="78" swimtime="00:00:56.99" resultid="3421" heatid="4645" lane="4" />
                <RESULT eventid="1074" points="130" swimtime="00:00:49.72" resultid="3422" heatid="4700" lane="2" entrytime="00:00:50.97" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucca" lastname="Diedrichs Santos" birthdate="2011-10-27" gender="M" nation="BRA" license="414417" swrid="5755372" athleteid="3451" externalid="414417" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="3452" heatid="4769" lane="4" />
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="3453" heatid="4829" lane="6" />
                <RESULT eventid="1213" status="DNS" swimtime="00:00:00.00" resultid="3454" heatid="4946" lane="4" />
                <RESULT eventid="1263" status="DNS" swimtime="00:00:00.00" resultid="3455" heatid="4992" lane="4" />
                <RESULT eventid="1329" status="DNS" swimtime="00:00:00.00" resultid="3457" heatid="5137" lane="5" />
                <RESULT eventid="10332" points="384" swimtime="00:00:27.72" resultid="10480" heatid="10347" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruna" lastname="Scalise Drapzichinski" birthdate="2012-03-07" gender="F" nation="BRA" license="378349" swrid="5603909" athleteid="3113" externalid="378349" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="382" swimtime="00:00:33.60" resultid="3114" heatid="4677" lane="6" entrytime="00:00:35.11" entrycourse="SCM" />
                <RESULT eventid="1077" points="290" swimtime="00:00:38.12" resultid="3115" heatid="4728" lane="1" entrytime="00:00:39.38" entrycourse="SCM" />
                <RESULT eventid="1129" points="431" swimtime="00:01:22.51" resultid="3116" heatid="4890" lane="4" entrytime="00:01:22.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="376" swimtime="00:03:06.44" resultid="3117" heatid="4923" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                    <SPLIT distance="100" swimtime="00:01:26.17" />
                    <SPLIT distance="150" swimtime="00:02:15.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="386" swimtime="00:00:31.47" resultid="3118" heatid="5103" lane="2" entrytime="00:00:30.55" entrycourse="SCM" />
                <RESULT eventid="1301" points="419" swimtime="00:00:37.91" resultid="3119" heatid="5051" lane="4" entrytime="00:00:37.39" entrycourse="SCM" />
                <RESULT eventid="4411" points="373" swimtime="00:00:33.86" resultid="5614" heatid="4681" lane="2" />
                <RESULT eventid="4413" points="375" swimtime="00:00:33.80" resultid="5636" heatid="4691" lane="4" />
                <RESULT eventid="4417" points="314" swimtime="00:00:37.14" resultid="5656" heatid="4732" lane="1" />
                <RESULT eventid="4419" points="318" swimtime="00:00:36.99" resultid="5680" heatid="4742" lane="4" />
                <RESULT eventid="5801" points="419" swimtime="00:00:37.89" resultid="10017" heatid="6069" lane="1" />
                <RESULT eventid="5804" points="384" swimtime="00:00:31.52" resultid="10056" heatid="6055" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Sprengel Betim" birthdate="2012-08-17" gender="F" nation="BRA" license="385011" swrid="5588922" athleteid="3348" externalid="385011" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="251" swimtime="00:00:38.60" resultid="3349" heatid="4669" lane="5" entrytime="00:00:38.75" entrycourse="SCM" />
                <RESULT eventid="1077" points="188" swimtime="00:00:44.07" resultid="3350" heatid="4711" lane="4" />
                <RESULT eventid="1179" points="256" swimtime="00:03:31.80" resultid="3351" heatid="4920" lane="1" />
                <RESULT eventid="1153" points="215" swimtime="00:01:30.17" resultid="3352" heatid="4900" lane="3" entrytime="00:01:42.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="265" swimtime="00:00:35.67" resultid="3353" heatid="5090" lane="6" entrytime="00:00:35.06" entrycourse="SCM" />
                <RESULT eventid="1301" points="223" swimtime="00:00:46.75" resultid="3354" heatid="5037" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Henrique Ballatka" birthdate="2013-08-26" gender="M" nation="BRA" license="405839" swrid="5697229" athleteid="3321" externalid="405839" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="41" swimtime="00:01:02.68" resultid="3322" heatid="4773" lane="6" />
                <RESULT eventid="1105" points="69" swimtime="00:00:53.87" resultid="3323" heatid="4833" lane="2" />
                <RESULT eventid="1273" points="91" swimtime="00:01:39.68" resultid="3324" heatid="5003" lane="5" entrytime="00:01:48.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.29" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida." eventid="1329" status="DSQ" swimtime="00:00:51.70" resultid="3326" heatid="5148" lane="6" entrytime="00:01:17.25" entrycourse="SCM" />
                <RESULT eventid="10332" points="92" swimtime="00:00:44.52" resultid="10472" heatid="10349" lane="6" entrytime="00:00:49.73" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Britto" birthdate="2012-10-04" gender="M" nation="BRA" license="378350" swrid="5588566" athleteid="3134" externalid="378350" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="228" swimtime="00:00:35.58" resultid="3135" heatid="4788" lane="3" entrytime="00:00:35.52" entrycourse="SCM" />
                <RESULT eventid="1105" points="223" swimtime="00:00:36.44" resultid="3136" heatid="4850" lane="1" entrytime="00:00:34.84" entrycourse="SCM" />
                <RESULT eventid="1203" points="225" swimtime="00:02:53.48" resultid="3137" heatid="4945" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                    <SPLIT distance="100" swimtime="00:01:24.98" />
                    <SPLIT distance="150" swimtime="00:02:10.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="217" swimtime="00:01:20.35" resultid="3138" heatid="4989" lane="1" entrytime="00:01:15.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="261" swimtime="00:00:31.51" resultid="3139" heatid="5222" lane="4" entrytime="00:00:31.01" entrycourse="SCM" />
                <RESULT eventid="1329" points="168" swimtime="00:00:45.18" resultid="3140" heatid="5157" lane="3" />
                <RESULT eventid="4423" points="227" swimtime="00:00:35.62" resultid="5702" heatid="4795" lane="4" />
                <RESULT eventid="4425" points="205" swimtime="00:00:36.86" resultid="5733" heatid="4805" lane="6" />
                <RESULT eventid="4429" points="214" swimtime="00:00:36.94" resultid="5752" heatid="4855" lane="2" />
                <RESULT eventid="4431" points="228" swimtime="00:00:36.18" resultid="5781" heatid="4865" lane="5" />
                <RESULT eventid="5807" points="177" swimtime="00:00:44.43" resultid="10131" heatid="6039" lane="5" />
                <RESULT eventid="5810" points="264" swimtime="00:00:31.39" resultid="10241" heatid="6023" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiggi" lastname="Frasson Abreu" birthdate="2014-07-16" gender="M" nation="BRA" license="411413" swrid="5077239" athleteid="3437" externalid="411413" level="MRGA">
              <RESULTS>
                <RESULT eventid="1089" points="28" swimtime="00:01:10.95" resultid="3438" heatid="4757" lane="3" entrytime="00:01:17.10" entrycourse="SCM" />
                <RESULT eventid="1102" points="37" swimtime="00:01:06.11" resultid="3439" heatid="4819" lane="5" entrytime="00:01:04.12" entrycourse="SCM" />
                <RESULT eventid="1213" points="55" swimtime="00:02:25.07" resultid="3440" heatid="4957" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="44" swimtime="00:02:06.90" resultid="3441" heatid="5012" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="43" swimtime="00:00:57.16" resultid="3442" heatid="5192" lane="2" entrytime="00:00:55.40" entrycourse="SCM" />
                <RESULT eventid="1326" points="54" swimtime="00:01:05.75" resultid="3443" heatid="5132" lane="3" entrytime="00:01:03.66" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Paes Schemiko" birthdate="2013-02-25" gender="F" nation="BRA" license="406918" swrid="5725995" athleteid="3375" externalid="406918" level="CLBO">
              <RESULTS>
                <RESULT comment="SW 8.2 - Braços não trazidos para frente simultaneamente sobre (em cima) a água." eventid="1064" status="DSQ" swimtime="00:00:38.45" resultid="3376" heatid="4668" lane="5" entrytime="00:00:40.01" entrycourse="SCM" />
                <RESULT eventid="1077" points="233" swimtime="00:00:40.98" resultid="3377" heatid="4718" lane="6" entrytime="00:00:41.48" entrycourse="SCM" />
                <RESULT eventid="1143" points="261" swimtime="00:02:52.56" resultid="3378" heatid="4893" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="265" swimtime="00:01:18.20" resultid="3379" heatid="4925" lane="3" />
                <RESULT eventid="1314" points="326" swimtime="00:00:33.31" resultid="3380" heatid="5090" lane="4" entrytime="00:00:33.76" entrycourse="SCM" />
                <RESULT eventid="1301" points="263" swimtime="00:00:44.27" resultid="3381" heatid="5041" lane="2" entrytime="00:00:47.05" entrycourse="SCM" />
                <RESULT eventid="5801" points="260" swimtime="00:00:44.40" resultid="10095" heatid="6066" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Schmeiske Ruivo" birthdate="2013-10-21" gender="F" nation="BRA" license="402006" swrid="5661354" athleteid="3309" externalid="402006" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="309" swimtime="00:00:36.03" resultid="3310" heatid="4674" lane="4" />
                <RESULT eventid="1077" points="274" swimtime="00:00:38.86" resultid="3311" heatid="4727" lane="4" entrytime="00:00:40.65" entrycourse="SCM" />
                <RESULT eventid="1129" points="323" swimtime="00:01:30.85" resultid="3312" heatid="4890" lane="2" entrytime="00:01:35.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="300" swimtime="00:03:20.92" resultid="3313" heatid="4923" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.96" />
                    <SPLIT distance="100" swimtime="00:01:36.42" />
                    <SPLIT distance="150" swimtime="00:02:28.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="302" swimtime="00:00:34.16" resultid="3314" heatid="5101" lane="4" entrytime="00:00:33.69" entrycourse="SCM" />
                <RESULT eventid="1301" points="339" swimtime="00:00:40.68" resultid="3315" heatid="5050" lane="6" entrytime="00:00:49.38" entrycourse="SCM" />
                <RESULT eventid="4411" points="316" swimtime="00:00:35.79" resultid="5607" heatid="4679" lane="1" />
                <RESULT eventid="4413" points="337" swimtime="00:00:35.01" resultid="5634" heatid="4690" lane="5" />
                <RESULT eventid="4417" points="272" swimtime="00:00:38.97" resultid="5651" heatid="4730" lane="2" />
                <RESULT eventid="4419" points="259" swimtime="00:00:39.57" resultid="5679" heatid="4741" lane="6" />
                <RESULT eventid="5801" points="317" swimtime="00:00:41.57" resultid="10011" heatid="6067" lane="1" />
                <RESULT eventid="5804" points="306" swimtime="00:00:34.01" resultid="10051" heatid="6053" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Ferreira Rais" birthdate="2007-07-04" gender="M" nation="BRA" license="398656" swrid="5697227" athleteid="3334" externalid="398656" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="415" swimtime="00:00:29.15" resultid="3335" heatid="4780" lane="5" entrytime="00:00:30.15" entrycourse="SCM" />
                <RESULT eventid="1105" points="265" swimtime="00:00:34.38" resultid="3336" heatid="4838" lane="6" entrytime="00:00:37.66" entrycourse="SCM" />
                <RESULT eventid="1237" points="296" swimtime="00:01:11.66" resultid="3337" heatid="4974" lane="6" entrytime="00:01:11.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="434" swimtime="00:00:59.22" resultid="3338" heatid="5009" lane="4" entrytime="00:01:01.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="219" swimtime="00:00:41.35" resultid="3340" heatid="5143" lane="6" />
                <RESULT eventid="10332" points="436" swimtime="00:00:26.57" resultid="10474" heatid="10358" lane="8" entrytime="00:00:26.77" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benicio" lastname="Garcia" birthdate="2011-09-09" gender="M" nation="BRA" license="378347" swrid="5603842" athleteid="3106" externalid="378347" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="207" swimtime="00:00:36.75" resultid="3107" heatid="4788" lane="1" entrytime="00:00:37.70" entrycourse="SCM" />
                <RESULT eventid="1105" points="227" swimtime="00:00:36.24" resultid="3108" heatid="4850" lane="6" entrytime="00:00:35.10" entrycourse="SCM" />
                <RESULT eventid="1249" points="238" swimtime="00:01:17.96" resultid="3109" heatid="4988" lane="4" entrytime="00:01:17.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1237" points="159" swimtime="00:01:28.08" resultid="3110" heatid="4976" lane="1" entrytime="00:01:38.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="281" swimtime="00:00:30.76" resultid="3111" heatid="5221" lane="5" entrytime="00:00:33.41" entrycourse="SCM" />
                <RESULT eventid="1329" points="163" swimtime="00:00:45.59" resultid="3112" heatid="5162" lane="5" entrytime="00:00:50.57" entrycourse="SCM" />
                <RESULT eventid="4429" points="267" swimtime="00:00:34.30" resultid="5760" heatid="4857" lane="4" />
                <RESULT eventid="4431" points="216" swimtime="00:00:36.83" resultid="5785" heatid="4866" lane="6" />
                <RESULT eventid="5810" points="272" swimtime="00:00:31.11" resultid="10249" heatid="6025" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dante" lastname="Gabriel Rossi" birthdate="2016-01-19" gender="M" nation="BRA" license="406928" swrid="5718627" athleteid="3403" externalid="406928" level="MRGA">
              <RESULTS>
                <RESULT eventid="1201" points="63" swimtime="00:00:55.56" resultid="3404" heatid="4941" lane="4" entrytime="00:01:00.59" entrycourse="SCM" />
                <RESULT eventid="1261" points="92" swimtime="00:00:44.61" resultid="3405" heatid="4991" lane="4" entrytime="00:00:46.06" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Gevaerd Verssutti Garcia" birthdate="2013-10-15" gender="F" nation="BRA" license="378404" swrid="5588723" athleteid="3239" externalid="378404" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="239" swimtime="00:00:39.27" resultid="3240" heatid="4673" lane="2" />
                <RESULT eventid="1077" points="255" swimtime="00:00:39.81" resultid="3241" heatid="4728" lane="6" entrytime="00:00:39.90" entrycourse="SCM" />
                <RESULT eventid="1119" status="DNS" swimtime="00:00:00.00" resultid="3242" heatid="4877" lane="4" />
                <RESULT eventid="1165" points="249" swimtime="00:01:27.20" resultid="3243" heatid="4917" lane="6" entrytime="00:01:29.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="259" swimtime="00:00:35.95" resultid="3244" heatid="5099" lane="3" entrytime="00:00:36.82" entrycourse="SCM" />
                <RESULT eventid="1301" points="167" swimtime="00:00:51.48" resultid="3245" heatid="5049" lane="2" entrytime="00:00:53.03" entrycourse="SCM" />
                <RESULT eventid="4411" points="248" swimtime="00:00:38.76" resultid="5611" heatid="4679" lane="5" />
                <RESULT eventid="4417" points="233" swimtime="00:00:41.01" resultid="5653" heatid="4730" lane="4" />
                <RESULT eventid="5801" points="159" swimtime="00:00:52.26" resultid="10016" heatid="6067" lane="6" />
                <RESULT eventid="5804" points="263" swimtime="00:00:35.78" resultid="10053" heatid="6053" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Berto" birthdate="2008-10-22" gender="M" nation="BRA" license="378342" swrid="5312223" athleteid="3183" externalid="378342" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="280" swimtime="00:00:33.24" resultid="3184" heatid="4789" lane="6" entrytime="00:00:35.22" entrycourse="SCM" />
                <RESULT eventid="1105" points="186" swimtime="00:00:38.71" resultid="3185" heatid="4847" lane="6" />
                <RESULT eventid="1213" points="331" swimtime="00:01:19.85" resultid="3186" heatid="4958" lane="3" entrytime="00:01:17.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="330" swimtime="00:02:53.85" resultid="3187" heatid="4995" lane="5" entrytime="00:02:43.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.73" />
                    <SPLIT distance="100" swimtime="00:01:23.17" />
                    <SPLIT distance="150" swimtime="00:02:07.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="296" swimtime="00:00:30.22" resultid="3188" heatid="5223" lane="1" entrytime="00:00:30.16" entrycourse="SCM" />
                <RESULT eventid="1329" points="331" swimtime="00:00:36.06" resultid="3189" heatid="5164" lane="4" entrytime="00:00:36.18" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Guidin Madureira" birthdate="2015-01-10" gender="M" nation="BRA" license="402116" swrid="5661347" athleteid="3316" externalid="402116" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="32" swimtime="00:01:08.04" resultid="3317" heatid="4751" lane="5" />
                <RESULT eventid="1102" points="71" swimtime="00:00:53.22" resultid="3318" heatid="4812" lane="3" entrytime="00:01:03.68" entrycourse="SCM" />
                <RESULT eventid="1326" points="52" swimtime="00:01:06.60" resultid="3320" heatid="5124" lane="7" />
                <RESULT eventid="10329" points="123" swimtime="00:00:40.49" resultid="10471" heatid="10342" lane="4" entrytime="00:00:43.45" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eloah" lastname="Juvedi Trindade" birthdate="2011-03-05" gender="F" nation="BRA" license="396829" swrid="5641768" athleteid="3281" externalid="396829" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="201" swimtime="00:00:41.59" resultid="3282" heatid="4674" lane="1" />
                <RESULT eventid="1077" points="230" swimtime="00:00:41.18" resultid="3283" heatid="4723" lane="5" />
                <RESULT eventid="1129" points="259" swimtime="00:01:37.73" resultid="3284" heatid="4890" lane="5" entrytime="00:01:36.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="232" swimtime="00:01:29.21" resultid="3285" heatid="4917" lane="1" entrytime="00:01:27.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="271" swimtime="00:00:35.40" resultid="3286" heatid="5102" lane="6" entrytime="00:00:33.38" entrycourse="SCM" />
                <RESULT eventid="1301" points="229" swimtime="00:00:46.31" resultid="3287" heatid="5048" lane="2" />
                <RESULT eventid="4411" points="195" swimtime="00:00:42.02" resultid="5621" heatid="4683" lane="3" />
                <RESULT eventid="4417" points="240" swimtime="00:00:40.63" resultid="5663" heatid="4734" lane="2" />
                <RESULT eventid="4419" points="248" swimtime="00:00:40.15" resultid="5685" heatid="4743" lane="6" />
                <RESULT eventid="5801" points="242" swimtime="00:00:45.48" resultid="10023" heatid="6071" lane="1" />
                <RESULT eventid="5804" points="268" swimtime="00:00:35.55" resultid="10062" heatid="6057" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Jupi Takaki" birthdate="2013-03-26" gender="F" nation="BRA" license="391845" swrid="5603861" athleteid="3260" externalid="391845" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="289" swimtime="00:00:36.85" resultid="3261" heatid="4676" lane="4" entrytime="00:00:36.53" entrycourse="SCM" />
                <RESULT eventid="1077" points="211" swimtime="00:00:42.39" resultid="3262" heatid="4723" lane="1" />
                <RESULT eventid="1153" points="236" swimtime="00:01:27.45" resultid="3263" heatid="4903" lane="6" entrytime="00:01:30.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="240" swimtime="00:01:20.76" resultid="3264" heatid="4937" lane="1" entrytime="00:01:24.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="263" swimtime="00:00:35.78" resultid="3265" heatid="5099" lane="4" entrytime="00:00:36.91" entrycourse="SCM" />
                <RESULT eventid="1301" points="144" swimtime="00:00:54.01" resultid="3266" heatid="5048" lane="3" />
                <RESULT eventid="4411" points="292" swimtime="00:00:36.73" resultid="5609" heatid="4679" lane="3" />
                <RESULT eventid="4417" points="227" swimtime="00:00:41.37" resultid="5654" heatid="4730" lane="5" />
                <RESULT eventid="5804" points="264" swimtime="00:00:35.74" resultid="10052" heatid="6053" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Drapzichinski" birthdate="2015-08-21" gender="M" nation="BRA" license="391848" swrid="5603890" athleteid="3267" externalid="391848" level="MRGA">
              <RESULTS>
                <RESULT eventid="1089" points="85" swimtime="00:00:49.33" resultid="3268" heatid="4757" lane="2" />
                <RESULT eventid="1102" points="108" swimtime="00:00:46.41" resultid="3269" heatid="4820" lane="4" entrytime="00:00:45.94" entrycourse="SCM" />
                <RESULT eventid="1249" points="97" swimtime="00:01:44.84" resultid="3270" heatid="4987" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="109" swimtime="00:01:33.69" resultid="3271" heatid="5013" lane="5" entrytime="00:01:38.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="129" swimtime="00:00:39.84" resultid="3272" heatid="5194" lane="2" entrytime="00:00:37.75" entrycourse="SCM" />
                <RESULT eventid="1326" points="78" swimtime="00:00:58.30" resultid="3273" heatid="5133" lane="5" entrytime="00:00:56.86" entrycourse="SCM" />
                <RESULT eventid="4421" points="109" swimtime="00:00:45.48" resultid="9024" heatid="9005" lane="6" />
                <RESULT eventid="4427" points="103" swimtime="00:00:47.15" resultid="9028" heatid="9007" lane="4" />
                <RESULT eventid="4445" points="84" swimtime="00:00:56.92" resultid="10113" heatid="6033" lane="3" />
                <RESULT eventid="4451" points="134" swimtime="00:00:39.33" resultid="10224" heatid="6017" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Manoel Forte" birthdate="2013-01-13" gender="M" nation="BRA" license="414859" swrid="5755340" athleteid="3464" externalid="414859" level="CLBO">
              <RESULTS>
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente., Na volta dos 25m." eventid="1092" status="DSQ" swimtime="00:01:03.27" resultid="3465" heatid="4771" lane="4" />
                <RESULT eventid="1105" points="90" swimtime="00:00:49.27" resultid="3466" heatid="4830" lane="5" />
                <RESULT eventid="1227" points="110" swimtime="00:03:26.98" resultid="3467" heatid="4964" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.18" />
                    <SPLIT distance="100" swimtime="00:01:38.16" />
                    <SPLIT distance="150" swimtime="00:02:33.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="103" swimtime="00:01:35.65" resultid="3468" heatid="4999" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" status="DNS" swimtime="00:00:00.00" resultid="3470" heatid="5146" lane="7" />
                <RESULT eventid="10332" status="DNS" swimtime="00:00:00.00" resultid="10481" heatid="10348" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Posser" birthdate="2013-02-07" gender="F" nation="BRA" license="378343" swrid="5603896" athleteid="3211" externalid="378343" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="196" swimtime="00:00:41.97" resultid="3212" heatid="4675" lane="2" entrytime="00:00:43.43" entrycourse="SCM" />
                <RESULT eventid="1077" points="139" swimtime="00:00:48.72" resultid="3213" heatid="4723" lane="6" />
                <RESULT eventid="1153" points="152" swimtime="00:01:41.22" resultid="3214" heatid="4902" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="212" swimtime="00:01:24.23" resultid="3215" heatid="4937" lane="5" entrytime="00:01:24.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="234" swimtime="00:00:37.17" resultid="3216" heatid="5098" lane="4" entrytime="00:00:42.80" entrycourse="SCM" />
                <RESULT eventid="1301" points="179" swimtime="00:00:50.28" resultid="3217" heatid="5047" lane="6" />
                <RESULT eventid="4411" points="191" swimtime="00:00:42.32" resultid="5612" heatid="4679" lane="6" />
                <RESULT eventid="5801" points="179" swimtime="00:00:50.26" resultid="10014" heatid="6067" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kauana" lastname="De Leal" birthdate="2016-02-20" gender="F" nation="BRA" license="417997" athleteid="3478" externalid="417997" level="MRGA">
              <RESULTS>
                <RESULT eventid="1177" points="33" swimtime="00:01:11.44" resultid="3479" heatid="4919" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marco" lastname="Manzotti Marchi" birthdate="2015-06-26" gender="M" nation="BRA" license="396849" swrid="5641769" athleteid="3288" externalid="396849" level="MRGA">
              <RESULTS>
                <RESULT eventid="1089" points="101" swimtime="00:00:46.68" resultid="3289" heatid="4759" lane="6" entrytime="00:00:52.83" entrycourse="SCM" />
                <RESULT eventid="1102" points="55" swimtime="00:00:58.10" resultid="3290" heatid="4819" lane="1" />
                <RESULT eventid="1237" points="74" swimtime="00:01:53.61" resultid="3291" heatid="4975" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="88" swimtime="00:01:40.57" resultid="3292" heatid="5012" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1285" points="94" swimtime="00:00:44.19" resultid="3293" heatid="5192" lane="5" />
                <RESULT eventid="1326" points="71" swimtime="00:01:00.13" resultid="3294" heatid="5132" lane="5" />
                <RESULT eventid="4421" points="96" swimtime="00:00:47.45" resultid="9022" heatid="9005" lane="4" />
                <RESULT eventid="4445" points="76" swimtime="00:00:58.74" resultid="10114" heatid="6033" lane="4" />
                <RESULT eventid="4451" points="94" swimtime="00:00:44.29" resultid="10227" heatid="6017" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Livia" lastname="Eloisa Silva" birthdate="2012-03-03" gender="F" nation="BRA" license="399725" swrid="5651341" athleteid="3302" externalid="399725" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="109" swimtime="00:00:50.99" resultid="3303" heatid="4674" lane="3" />
                <RESULT eventid="1077" points="148" swimtime="00:00:47.70" resultid="3304" heatid="4725" lane="2" entrytime="00:00:50.69" entrycourse="SCM" />
                <RESULT eventid="1165" points="152" swimtime="00:01:42.80" resultid="3305" heatid="4916" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="113" swimtime="00:01:43.89" resultid="3306" heatid="4934" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="114" swimtime="00:00:47.16" resultid="3307" heatid="5098" lane="2" entrytime="00:00:45.25" entrycourse="SCM" />
                <RESULT eventid="1301" points="37" swimtime="00:01:24.93" resultid="3308" heatid="5047" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Rezende" birthdate="2012-01-23" gender="F" nation="BRA" license="370669" swrid="5603899" athleteid="3232" externalid="370669" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="109" swimtime="00:00:50.97" resultid="3233" heatid="4674" lane="6" />
                <RESULT eventid="1077" points="196" swimtime="00:00:43.41" resultid="3234" heatid="4725" lane="3" entrytime="00:00:46.31" entrycourse="SCM" />
                <RESULT eventid="1119" points="212" swimtime="00:03:19.46" resultid="3235" heatid="4877" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.71" />
                    <SPLIT distance="100" swimtime="00:01:37.26" />
                    <SPLIT distance="150" swimtime="00:02:28.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="210" swimtime="00:01:24.47" resultid="3236" heatid="4938" lane="1" entrytime="00:01:18.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="221" swimtime="00:00:37.92" resultid="3237" heatid="5100" lane="3" entrytime="00:00:34.83" entrycourse="SCM" />
                <RESULT eventid="1301" points="209" swimtime="00:00:47.73" resultid="3238" heatid="5049" lane="3" entrytime="00:00:50.89" entrycourse="SCM" />
                <RESULT eventid="4417" status="DNS" swimtime="00:00:00.00" resultid="5660" heatid="4732" lane="5" />
                <RESULT eventid="5801" points="204" swimtime="00:00:48.16" resultid="10022" heatid="6069" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Zanatta Duda" birthdate="2013-08-28" gender="F" nation="BRA" license="406914" swrid="5717306" athleteid="3362" externalid="406914" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="96" swimtime="00:00:53.18" resultid="3363" heatid="4663" lane="3" />
                <RESULT eventid="1077" points="169" swimtime="00:00:45.65" resultid="3364" heatid="4715" lane="4" entrytime="00:00:46.45" entrycourse="SCM" />
                <RESULT eventid="1189" points="176" swimtime="00:01:29.55" resultid="3365" heatid="4928" lane="6" entrytime="00:01:33.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="199" swimtime="00:00:39.21" resultid="3366" heatid="5086" lane="1" entrytime="00:00:40.92" entrycourse="SCM" />
                <RESULT eventid="1301" points="86" swimtime="00:01:04.23" resultid="3367" heatid="5037" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Guilherme Ballatka" birthdate="2007-06-24" gender="M" nation="BRA" license="398616" swrid="5697228" athleteid="3327" externalid="398616" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="324" swimtime="00:00:31.66" resultid="3328" heatid="4764" lane="1" />
                <RESULT eventid="1105" points="418" swimtime="00:00:29.57" resultid="3329" heatid="4841" lane="3" entrytime="00:00:28.76" entrycourse="SCM" />
                <RESULT eventid="1203" points="412" swimtime="00:02:21.93" resultid="3330" heatid="4943" lane="3" entrytime="00:02:17.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.31" />
                    <SPLIT distance="100" swimtime="00:01:07.07" />
                    <SPLIT distance="150" swimtime="00:01:44.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="435" swimtime="00:01:03.74" resultid="3331" heatid="4986" lane="3" entrytime="00:01:03.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="373" swimtime="00:00:34.64" resultid="3333" heatid="5140" lane="3" />
                <RESULT eventid="4429" points="441" swimtime="00:00:29.04" resultid="5591" heatid="4862" lane="1" />
                <RESULT eventid="4431" points="390" swimtime="00:00:30.25" resultid="5597" heatid="4869" lane="1" />
                <RESULT eventid="5807" points="368" swimtime="00:00:34.81" resultid="10303" heatid="6046" lane="5" />
                <RESULT eventid="10332" points="476" swimtime="00:00:25.81" resultid="10473" heatid="10360" lane="6" entrytime="00:00:25.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernanda" lastname="Camillo Sabim" birthdate="2010-08-02" gender="F" nation="BRA" license="406931" swrid="5723021" athleteid="3406" externalid="406931" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="193" swimtime="00:00:42.16" resultid="3407" heatid="4660" lane="2" />
                <RESULT eventid="1077" points="265" swimtime="00:00:39.29" resultid="3408" heatid="4714" lane="6" />
                <RESULT eventid="1129" points="298" swimtime="00:01:33.34" resultid="3409" heatid="4884" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="322" swimtime="00:03:16.26" resultid="3410" heatid="4922" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.05" />
                    <SPLIT distance="100" swimtime="00:01:33.58" />
                    <SPLIT distance="150" swimtime="00:02:25.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="310" swimtime="00:00:33.87" resultid="3411" heatid="5085" lane="7" />
                <RESULT eventid="1301" points="321" swimtime="00:00:41.43" resultid="3412" heatid="5032" lane="3" />
                <RESULT eventid="4417" points="282" swimtime="00:00:38.49" resultid="5440" heatid="4735" lane="5" />
                <RESULT eventid="5801" points="327" swimtime="00:00:41.17" resultid="10107" heatid="6072" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Schneider Yazbek" birthdate="2013-03-07" gender="F" nation="BRA" license="378329" swrid="5588907" athleteid="3274" externalid="378329" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="288" swimtime="00:00:36.89" resultid="3275" heatid="4660" lane="3" />
                <RESULT eventid="1077" points="253" swimtime="00:00:39.90" resultid="3276" heatid="4717" lane="5" entrytime="00:00:41.99" entrycourse="SCM" />
                <RESULT eventid="1153" points="247" swimtime="00:01:26.05" resultid="3277" heatid="4901" lane="6" entrytime="00:01:33.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="411" swimtime="00:02:28.35" resultid="3278" heatid="4895" lane="2" entrytime="00:02:35.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                    <SPLIT distance="100" swimtime="00:01:12.73" />
                    <SPLIT distance="150" swimtime="00:01:51.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="358" swimtime="00:00:32.28" resultid="3279" heatid="5092" lane="2" entrytime="00:00:33.21" entrycourse="SCM" />
                <RESULT eventid="1301" points="230" swimtime="00:00:46.28" resultid="3280" heatid="5040" lane="4" entrytime="00:00:48.55" entrycourse="SCM" />
                <RESULT eventid="4411" points="318" swimtime="00:00:35.70" resultid="5385" heatid="4678" lane="5" />
                <RESULT eventid="4417" points="254" swimtime="00:00:39.86" resultid="5413" heatid="4729" lane="6" />
                <RESULT eventid="5804" points="372" swimtime="00:00:31.87" resultid="10188" heatid="6052" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Ognibeni Paupitz" birthdate="2014-08-08" gender="F" nation="BRA" license="406923" swrid="5718889" athleteid="3389" externalid="406923" level="MRGA">
              <RESULTS>
                <RESULT eventid="1061" points="71" swimtime="00:00:58.81" resultid="3390" heatid="4653" lane="6" />
                <RESULT eventid="1074" points="68" swimtime="00:01:01.85" resultid="3391" heatid="4704" lane="6" />
                <RESULT eventid="1129" points="112" swimtime="00:02:09.18" resultid="3392" heatid="4888" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="85" swimtime="00:01:54.21" resultid="3393" heatid="4934" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="125" swimtime="00:00:56.67" resultid="3394" heatid="5028" lane="5" entrytime="00:00:55.61" entrycourse="SCM" />
                <RESULT eventid="1311" points="132" swimtime="00:00:45.03" resultid="3395" heatid="5079" lane="6" entrytime="00:00:43.36" entrycourse="SCM" />
                <RESULT eventid="4433" points="130" swimtime="00:00:55.93" resultid="10009" heatid="6065" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Kuhnen Consalter" birthdate="2014-04-25" gender="F" nation="BRA" license="415372" swrid="5755357" athleteid="3471" externalid="415372" level="MRGA">
              <RESULTS>
                <RESULT eventid="1061" status="DNS" swimtime="00:00:00.00" resultid="3472" heatid="4654" lane="4" entrytime="00:00:45.73" entrycourse="SCM" />
                <RESULT eventid="1074" status="DNS" swimtime="00:00:00.00" resultid="3473" heatid="4703" lane="2" />
                <RESULT eventid="1129" status="DNS" swimtime="00:00:00.00" resultid="3474" heatid="4888" lane="6" />
                <RESULT eventid="1189" status="DNS" swimtime="00:00:00.00" resultid="3475" heatid="4935" lane="1" />
                <RESULT eventid="1298" status="DNS" swimtime="00:00:00.00" resultid="3476" heatid="5026" lane="4" />
                <RESULT eventid="1311" status="DNS" swimtime="00:00:00.00" resultid="3477" heatid="5079" lane="2" entrytime="00:00:38.79" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eloah" lastname="Frasson" birthdate="2012-06-14" gender="F" nation="BRA" license="378338" swrid="5577016" athleteid="3204" externalid="378338" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="224" swimtime="00:00:40.14" resultid="3205" heatid="4673" lane="3" />
                <RESULT eventid="1077" points="145" swimtime="00:00:48.05" resultid="3206" heatid="4723" lane="2" />
                <RESULT eventid="1129" points="299" swimtime="00:01:33.18" resultid="3207" heatid="4890" lane="6" entrytime="00:01:37.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="260" swimtime="00:01:18.64" resultid="3208" heatid="4937" lane="4" entrytime="00:01:22.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="237" swimtime="00:00:37.02" resultid="3209" heatid="5100" lane="1" entrytime="00:00:36.19" entrycourse="SCM" />
                <RESULT eventid="1301" points="308" swimtime="00:00:42.00" resultid="3210" heatid="5051" lane="6" entrytime="00:00:41.90" entrycourse="SCM" />
                <RESULT eventid="4411" points="224" swimtime="00:00:40.10" resultid="5618" heatid="4681" lane="6" />
                <RESULT eventid="5801" points="306" swimtime="00:00:42.08" resultid="10018" heatid="6069" lane="2" />
                <RESULT eventid="5804" points="269" swimtime="00:00:35.49" resultid="10061" heatid="6055" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aline" lastname="Hirano" birthdate="2007-11-13" gender="F" nation="BRA" license="358898" swrid="5622283" athleteid="3355" externalid="358898" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="331" swimtime="00:00:35.23" resultid="3356" heatid="4663" lane="2" />
                <RESULT eventid="1077" points="295" swimtime="00:00:37.90" resultid="3357" heatid="4711" lane="2" />
                <RESULT eventid="1179" points="276" swimtime="00:03:26.51" resultid="3358" heatid="4922" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.05" />
                    <SPLIT distance="100" swimtime="00:01:37.47" />
                    <SPLIT distance="150" swimtime="00:02:32.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="260" swimtime="00:01:24.63" resultid="3359" heatid="4899" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="390" swimtime="00:00:31.37" resultid="3360" heatid="5094" lane="2" entrytime="00:00:30.96" entrycourse="SCM" />
                <RESULT eventid="1301" status="DNS" swimtime="00:00:00.00" resultid="3361" heatid="5038" lane="5" />
                <RESULT eventid="4411" points="342" swimtime="00:00:34.86" resultid="5347" heatid="4688" lane="4" />
                <RESULT eventid="4417" points="376" swimtime="00:00:34.98" resultid="5458" heatid="4739" lane="5" />
                <RESULT eventid="4419" points="307" swimtime="00:00:37.40" resultid="5462" heatid="4746" lane="3" />
                <RESULT eventid="5804" points="385" swimtime="00:00:31.50" resultid="10216" heatid="6062" lane="5" />
                <RESULT eventid="4413" points="228" swimtime="00:00:39.87" resultid="10322" heatid="4695" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Ribeiro Melo" birthdate="2011-07-01" gender="F" nation="BRA" license="390923" swrid="5602577" athleteid="3148" externalid="390923" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="336" swimtime="00:00:35.04" resultid="3149" heatid="4670" lane="1" entrytime="00:00:37.28" entrycourse="SCM" />
                <RESULT eventid="1077" points="313" swimtime="00:00:37.15" resultid="3150" heatid="4720" lane="1" entrytime="00:00:38.48" entrycourse="SCM" />
                <RESULT eventid="1129" points="309" swimtime="00:01:32.17" resultid="3151" heatid="4885" lane="4" entrytime="00:01:35.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="271" swimtime="00:01:24.73" resultid="3152" heatid="4911" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="386" swimtime="00:00:31.49" resultid="3153" heatid="5096" lane="1" entrytime="00:00:30.60" entrycourse="SCM" />
                <RESULT eventid="1301" points="295" swimtime="00:00:42.59" resultid="3154" heatid="5042" lane="8" entrytime="00:00:42.69" entrycourse="SCM" />
                <RESULT eventid="4411" points="336" swimtime="00:00:35.04" resultid="5354" heatid="4682" lane="2" />
                <RESULT eventid="4413" points="262" swimtime="00:00:38.08" resultid="5360" heatid="4692" lane="2" />
                <RESULT eventid="5804" points="408" swimtime="00:00:30.90" resultid="10202" heatid="6056" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Valentina Gozaga" birthdate="2014-06-28" gender="F" nation="BRA" license="385709" swrid="5603924" athleteid="3253" externalid="385709" level="MRGA">
              <RESULTS>
                <RESULT eventid="1061" points="63" swimtime="00:01:01.14" resultid="3254" heatid="4652" lane="2" />
                <RESULT eventid="1074" points="147" swimtime="00:00:47.77" resultid="3255" heatid="4705" lane="2" entrytime="00:00:47.42" entrycourse="SCM" />
                <RESULT eventid="1129" points="145" swimtime="00:01:58.48" resultid="3256" heatid="4889" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="115" swimtime="00:01:52.74" resultid="3257" heatid="4916" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="129" swimtime="00:00:56.07" resultid="3258" heatid="5028" lane="4" entrytime="00:00:53.76" entrycourse="SCM" />
                <RESULT eventid="1311" points="187" swimtime="00:00:40.06" resultid="3259" heatid="5079" lane="5" entrytime="00:00:39.26" entrycourse="SCM" />
                <RESULT eventid="4415" points="136" swimtime="00:00:49.09" resultid="9021" heatid="9004" lane="6" />
                <RESULT eventid="4433" points="148" swimtime="00:00:53.53" resultid="10008" heatid="6065" lane="4" />
                <RESULT eventid="4439" points="196" swimtime="00:00:39.41" resultid="10046" heatid="6051" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Laura Oliveira" birthdate="2014-05-19" gender="F" nation="BRA" license="414179" swrid="5336453" athleteid="3444" externalid="414179" level="MRGA">
              <RESULTS>
                <RESULT eventid="1061" points="82" swimtime="00:00:55.96" resultid="3445" heatid="4654" lane="6" entrytime="00:01:01.46" entrycourse="SCM" />
                <RESULT eventid="1074" points="87" swimtime="00:00:56.89" resultid="3446" heatid="4704" lane="3" entrytime="00:00:56.86" entrycourse="SCM" />
                <RESULT eventid="1165" points="91" swimtime="00:02:02.02" resultid="3447" heatid="4915" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="135" swimtime="00:01:37.79" resultid="3448" heatid="4936" lane="1" entrytime="00:01:50.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="41" swimtime="00:01:22.17" resultid="3449" heatid="5026" lane="2" />
                <RESULT eventid="1311" points="151" swimtime="00:00:43.03" resultid="3450" heatid="5078" lane="5" entrytime="00:00:46.77" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1115" points="249" swimtime="00:04:44.96" resultid="3494" heatid="5251" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                    <SPLIT distance="100" swimtime="00:01:20.57" />
                    <SPLIT distance="150" swimtime="00:01:50.41" />
                    <SPLIT distance="200" swimtime="00:02:28.42" />
                    <SPLIT distance="250" swimtime="00:03:04.70" />
                    <SPLIT distance="300" swimtime="00:03:34.91" />
                    <SPLIT distance="350" swimtime="00:04:07.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3197" number="1" />
                    <RELAYPOSITION athleteid="3267" number="2" />
                    <RELAYPOSITION athleteid="3155" number="3" />
                    <RELAYPOSITION athleteid="3341" number="4" />
                    <RELAYPOSITION athleteid="3134" number="5" />
                    <RELAYPOSITION athleteid="3162" number="6" />
                    <RELAYPOSITION athleteid="3092" number="7" />
                    <RELAYPOSITION athleteid="3430" number="8" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1339" points="260" swimtime="00:04:16.04" resultid="3495" heatid="5252" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.83" />
                    <SPLIT distance="100" swimtime="00:01:06.80" />
                    <SPLIT distance="150" swimtime="00:01:44.22" />
                    <SPLIT distance="200" swimtime="00:02:23.62" />
                    <SPLIT distance="250" swimtime="00:02:50.90" />
                    <SPLIT distance="300" swimtime="00:03:22.57" />
                    <SPLIT distance="350" swimtime="00:03:49.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3197" number="1" />
                    <RELAYPOSITION athleteid="3341" number="2" />
                    <RELAYPOSITION athleteid="3430" number="3" />
                    <RELAYPOSITION athleteid="3267" number="4" />
                    <RELAYPOSITION athleteid="3092" number="5" />
                    <RELAYPOSITION athleteid="3134" number="6" />
                    <RELAYPOSITION athleteid="3162" number="7" />
                    <RELAYPOSITION athleteid="3155" number="8" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="FÁBRICA DE NADADORES &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1115" points="134" status="EXH" swimtime="00:05:49.81" resultid="3498" heatid="4871" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                    <SPLIT distance="100" swimtime="00:01:16.89" />
                    <SPLIT distance="150" swimtime="00:02:19.52" />
                    <SPLIT distance="200" swimtime="00:02:49.15" />
                    <SPLIT distance="250" swimtime="00:03:34.78" />
                    <SPLIT distance="300" swimtime="00:04:21.45" />
                    <SPLIT distance="350" swimtime="00:05:14.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3464" number="1" />
                    <RELAYPOSITION athleteid="3368" number="2" />
                    <RELAYPOSITION athleteid="3327" number="3" />
                    <RELAYPOSITION athleteid="3382" number="4" />
                    <RELAYPOSITION athleteid="3334" number="5" />
                    <RELAYPOSITION athleteid="3480" number="6" />
                    <RELAYPOSITION athleteid="3321" number="7" />
                    <RELAYPOSITION athleteid="3316" number="8" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1339" points="183" status="EXH" swimtime="00:04:48.11" resultid="3499" heatid="5246" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.05" />
                    <SPLIT distance="100" swimtime="00:01:00.12" />
                    <SPLIT distance="150" swimtime="00:01:41.80" />
                    <SPLIT distance="200" swimtime="00:02:26.92" />
                    <SPLIT distance="250" swimtime="00:03:04.09" />
                    <SPLIT distance="300" swimtime="00:03:35.73" />
                    <SPLIT distance="350" swimtime="00:04:21.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" />
                    <RELAYPOSITION number="2" reactiontime="0" />
                    <RELAYPOSITION number="3" reactiontime="0" />
                    <RELAYPOSITION number="4" reactiontime="0" />
                    <RELAYPOSITION number="5" reactiontime="0" />
                    <RELAYPOSITION number="6" reactiontime="0" />
                    <RELAYPOSITION number="7" reactiontime="0" />
                    <RELAYPOSITION number="8" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="FÁBRICA DE NADADORES &quot;C&quot;" number="3">
              <RESULTS>
                <RESULT eventid="1115" points="136" status="EXH" swimtime="00:05:48.59" resultid="5796" heatid="5251" lane="6" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.93" />
                    <SPLIT distance="100" swimtime="00:01:47.11" />
                    <SPLIT distance="150" swimtime="00:02:41.49" />
                    <SPLIT distance="200" swimtime="00:03:21.84" />
                    <SPLIT distance="250" swimtime="00:03:50.85" />
                    <SPLIT distance="300" swimtime="00:04:25.83" />
                    <SPLIT distance="350" swimtime="00:05:10.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3288" number="1" />
                    <RELAYPOSITION athleteid="3396" number="2" />
                    <RELAYPOSITION athleteid="3437" number="3" />
                    <RELAYPOSITION athleteid="3218" number="4" />
                    <RELAYPOSITION athleteid="3190" number="5" />
                    <RELAYPOSITION athleteid="3106" number="6" />
                    <RELAYPOSITION athleteid="3120" number="7" />
                    <RELAYPOSITION athleteid="3183" number="8" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1339" points="167" status="EXH" swimtime="00:04:56.70" resultid="10110" heatid="5252" lane="6" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                    <SPLIT distance="100" swimtime="00:01:12.86" />
                    <SPLIT distance="150" swimtime="00:02:07.63" />
                    <SPLIT distance="200" swimtime="00:02:39.29" />
                    <SPLIT distance="250" swimtime="00:03:23.11" />
                    <SPLIT distance="300" swimtime="00:03:55.19" />
                    <SPLIT distance="350" swimtime="00:04:26.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3190" number="1" />
                    <RELAYPOSITION athleteid="3288" number="2" />
                    <RELAYPOSITION athleteid="3437" number="3" />
                    <RELAYPOSITION athleteid="3169" number="4" />
                    <RELAYPOSITION athleteid="3396" number="5" />
                    <RELAYPOSITION athleteid="3218" number="6" />
                    <RELAYPOSITION athleteid="3106" number="7" />
                    <RELAYPOSITION athleteid="3183" number="8" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT comment="SW 10.12 - Os pés perderam contato com a plataforma de partida antes que o colega de equipe anterior tocasse a borda.  (Horário: 11:20)" eventid="1087" status="DSQ" swimtime="00:06:35.79" resultid="3492" heatid="5247" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.38" />
                    <SPLIT distance="100" swimtime="00:02:00.14" />
                    <SPLIT distance="150" swimtime="00:02:34.35" />
                    <SPLIT distance="200" swimtime="00:03:18.85" />
                    <SPLIT distance="250" swimtime="00:03:58.61" />
                    <SPLIT distance="300" swimtime="00:04:55.67" />
                    <SPLIT distance="350" swimtime="00:05:52.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3444" number="1" />
                    <RELAYPOSITION athleteid="3478" number="2" />
                    <RELAYPOSITION athleteid="3141" number="3" />
                    <RELAYPOSITION athleteid="3127" number="4" />
                    <RELAYPOSITION athleteid="3253" number="5" />
                    <RELAYPOSITION athleteid="3485" number="6" />
                    <RELAYPOSITION athleteid="3389" number="7" status="DSQ" />
                    <RELAYPOSITION athleteid="3204" number="8" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1324" points="276" swimtime="00:04:43.96" resultid="3493" heatid="5249" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.64" />
                    <SPLIT distance="100" swimtime="00:01:21.50" />
                    <SPLIT distance="150" swimtime="00:01:54.77" />
                    <SPLIT distance="200" swimtime="00:02:31.62" />
                    <SPLIT distance="250" swimtime="00:03:06.69" />
                    <SPLIT distance="300" swimtime="00:03:38.09" />
                    <SPLIT distance="350" swimtime="00:04:09.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3295" number="1" />
                    <RELAYPOSITION athleteid="3309" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3225" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3281" number="4" reactiontime="0" />
                    <RELAYPOSITION athleteid="3246" number="5" reactiontime="0" />
                    <RELAYPOSITION athleteid="3141" number="6" reactiontime="0" />
                    <RELAYPOSITION athleteid="3113" number="7" reactiontime="0" />
                    <RELAYPOSITION athleteid="3239" number="8" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="FÁBRICA DE NADADORES &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1087" points="277" swimtime="00:05:13.80" resultid="3496" heatid="5247" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.08" />
                    <SPLIT distance="100" swimtime="00:01:27.28" />
                    <SPLIT distance="150" swimtime="00:02:08.27" />
                    <SPLIT distance="200" swimtime="00:02:45.75" />
                    <SPLIT distance="250" swimtime="00:03:24.48" />
                    <SPLIT distance="300" swimtime="00:04:00.92" />
                    <SPLIT distance="350" swimtime="00:04:37.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3295" number="1" />
                    <RELAYPOSITION athleteid="3225" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3309" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3260" number="4" reactiontime="0" />
                    <RELAYPOSITION athleteid="3113" number="5" reactiontime="0" />
                    <RELAYPOSITION athleteid="3176" number="6" reactiontime="0" />
                    <RELAYPOSITION athleteid="3204" number="7" reactiontime="0" />
                    <RELAYPOSITION athleteid="3232" number="8" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1324" points="169" swimtime="00:05:34.26" resultid="3497" heatid="5249" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                    <SPLIT distance="100" swimtime="00:01:11.43" />
                    <SPLIT distance="150" swimtime="00:02:20.11" />
                    <SPLIT distance="200" swimtime="00:03:01.11" />
                    <SPLIT distance="250" swimtime="00:03:37.32" />
                    <SPLIT distance="300" swimtime="00:04:14.22" />
                    <SPLIT distance="350" swimtime="00:04:58.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3204" number="1" />
                    <RELAYPOSITION athleteid="3232" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3478" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3253" number="4" reactiontime="0" />
                    <RELAYPOSITION athleteid="3260" number="5" reactiontime="0" />
                    <RELAYPOSITION athleteid="3413" number="6" reactiontime="0" />
                    <RELAYPOSITION athleteid="3302" number="7" reactiontime="0" />
                    <RELAYPOSITION athleteid="3211" number="8" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="263" nation="BRA" region="PR" clubid="2182" swrid="75436" name="Clube Curitibano" shortname="Curitibano">
          <ATHLETES>
            <ATHLETE firstname="Lorenzo" lastname="Kraemer Geremia" birthdate="2013-08-16" gender="M" nation="BRA" license="377041" swrid="5588762" athleteid="2524" externalid="377041" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="218" swimtime="00:00:36.10" resultid="2525" heatid="4775" lane="3" entrytime="00:00:40.73" entrycourse="SCM" />
                <RESULT eventid="1105" points="227" swimtime="00:00:36.24" resultid="2526" heatid="4839" lane="1" entrytime="00:00:36.36" entrycourse="SCM" />
                <RESULT eventid="1203" points="230" swimtime="00:02:52.26" resultid="2527" heatid="4942" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.37" />
                    <SPLIT distance="100" swimtime="00:01:24.46" />
                    <SPLIT distance="150" swimtime="00:02:10.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="234" swimtime="00:01:18.36" resultid="2528" heatid="4985" lane="4" entrytime="00:01:22.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="183" swimtime="00:00:43.87" resultid="2530" heatid="5150" lane="4" entrytime="00:00:47.05" entrycourse="SCM" />
                <RESULT eventid="4423" points="192" swimtime="00:00:37.68" resultid="5483" heatid="4792" lane="3" />
                <RESULT eventid="4429" points="215" swimtime="00:00:36.89" resultid="5512" heatid="4852" lane="2" />
                <RESULT eventid="4431" points="225" swimtime="00:00:36.32" resultid="5518" heatid="4864" lane="2" />
                <RESULT eventid="5807" points="179" swimtime="00:00:44.22" resultid="10267" heatid="6036" lane="2" />
                <RESULT eventid="10332" points="265" swimtime="00:00:31.35" resultid="10427" heatid="10354" lane="2" entrytime="00:00:31.82" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Spadari Soso" birthdate="2012-12-28" gender="F" nation="BRA" license="377313" swrid="5588921" athleteid="2942" externalid="377313" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="280" swimtime="00:00:37.25" resultid="2943" heatid="4667" lane="1" entrytime="00:00:44.62" entrycourse="SCM" />
                <RESULT eventid="1077" points="245" swimtime="00:00:40.31" resultid="2944" heatid="4718" lane="3" entrytime="00:00:40.12" entrycourse="SCM" />
                <RESULT eventid="1143" points="414" swimtime="00:02:27.90" resultid="2945" heatid="4895" lane="6" entrytime="00:02:52.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.86" />
                    <SPLIT distance="100" swimtime="00:01:13.43" />
                    <SPLIT distance="150" swimtime="00:01:51.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="414" swimtime="00:01:07.41" resultid="2946" heatid="4931" lane="2" entrytime="00:01:10.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="383" swimtime="00:00:31.57" resultid="2947" heatid="5093" lane="4" entrytime="00:00:31.68" entrycourse="SCM" />
                <RESULT eventid="1301" points="310" swimtime="00:00:41.90" resultid="2948" heatid="5044" lane="8" entrytime="00:00:42.16" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Presiazniuk" birthdate="2010-10-14" gender="M" nation="BRA" license="356353" swrid="5600237" athleteid="2211" externalid="356353" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="256" swimtime="00:00:34.21" resultid="2212" heatid="4767" lane="2" />
                <RESULT eventid="1105" points="295" swimtime="00:00:33.20" resultid="2213" heatid="4840" lane="4" entrytime="00:00:31.92" entrycourse="SCM" />
                <RESULT eventid="1213" points="254" swimtime="00:01:27.22" resultid="2214" heatid="4949" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1237" points="248" swimtime="00:01:16.01" resultid="2215" heatid="4971" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="196" swimtime="00:00:42.88" resultid="2217" heatid="5142" lane="1" />
                <RESULT eventid="4429" points="302" swimtime="00:00:32.94" resultid="5578" heatid="4858" lane="3" />
                <RESULT eventid="4431" points="267" swimtime="00:00:34.31" resultid="5584" heatid="4867" lane="3" />
                <RESULT eventid="10332" points="375" swimtime="00:00:27.95" resultid="10402" heatid="10346" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernanda" lastname="Toscani Kim" birthdate="2013-02-15" gender="F" nation="BRA" license="372683" swrid="5588939" athleteid="2440" externalid="372683" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="281" swimtime="00:00:37.20" resultid="2441" heatid="4669" lane="3" entrytime="00:00:38.17" entrycourse="SCM" />
                <RESULT eventid="1077" points="232" swimtime="00:00:41.09" resultid="2442" heatid="4713" lane="6" />
                <RESULT eventid="1129" points="325" swimtime="00:01:30.62" resultid="2443" heatid="4886" lane="6" entrytime="00:01:31.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="313" swimtime="00:03:18.16" resultid="2444" heatid="4921" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.09" />
                    <SPLIT distance="100" swimtime="00:01:34.10" />
                    <SPLIT distance="150" swimtime="00:02:26.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="311" swimtime="00:00:33.81" resultid="2445" heatid="5089" lane="1" entrytime="00:00:35.39" entrycourse="SCM" />
                <RESULT eventid="1301" points="311" swimtime="00:00:41.83" resultid="2446" heatid="5042" lane="4" entrytime="00:00:43.14" entrycourse="SCM" />
                <RESULT eventid="4411" points="274" swimtime="00:00:37.50" resultid="5386" heatid="4678" lane="6" />
                <RESULT eventid="5801" points="305" swimtime="00:00:42.12" resultid="10094" heatid="6066" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Francia Soares" birthdate="2014-06-01" gender="F" nation="BRA" license="391011" swrid="5602540" athleteid="2636" externalid="391011" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" status="DNS" swimtime="00:00:00.00" resultid="2637" heatid="4647" lane="3" entrytime="00:01:06.21" entrycourse="SCM" />
                <RESULT eventid="1074" status="DNS" swimtime="00:00:00.00" resultid="2638" heatid="4699" lane="4" entrytime="00:00:53.98" entrycourse="SCM" />
                <RESULT eventid="1129" status="DNS" swimtime="00:00:00.00" resultid="2639" heatid="4883" lane="5" />
                <RESULT eventid="1189" status="DNS" swimtime="00:00:00.00" resultid="2640" heatid="4924" lane="2" />
                <RESULT eventid="1298" status="DNS" swimtime="00:00:00.00" resultid="2641" heatid="5020" lane="3" />
                <RESULT eventid="1311" status="DNS" swimtime="00:00:00.00" resultid="2642" heatid="5073" lane="5" entrytime="00:00:44.34" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Guimaraes Mesquita" birthdate="2013-12-30" gender="F" nation="BRA" license="391027" swrid="5602544" athleteid="2711" externalid="391027" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="93" swimtime="00:00:53.62" resultid="2712" heatid="4664" lane="2" />
                <RESULT eventid="1077" points="122" swimtime="00:00:50.80" resultid="2713" heatid="4709" lane="6" />
                <RESULT eventid="1129" points="172" swimtime="00:01:52.01" resultid="2714" heatid="4885" lane="1" entrytime="00:01:50.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="203" swimtime="00:03:48.84" resultid="2715" heatid="4920" lane="3" />
                <RESULT eventid="1314" points="209" swimtime="00:00:38.61" resultid="2716" heatid="5086" lane="5" entrytime="00:00:39.85" entrycourse="SCM" />
                <RESULT eventid="1301" points="185" swimtime="00:00:49.73" resultid="2717" heatid="5038" lane="8" entrytime="00:00:58.22" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Wolf Macedo" birthdate="2012-01-27" gender="F" nation="BRA" license="369277" swrid="5602592" athleteid="2384" externalid="369277" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="420" swimtime="00:00:32.54" resultid="2385" heatid="4671" lane="2" entrytime="00:00:33.20" entrycourse="SCM" />
                <RESULT eventid="1077" points="307" swimtime="00:00:37.41" resultid="2386" heatid="4719" lane="3" entrytime="00:00:38.96" entrycourse="SCM" />
                <RESULT eventid="1129" points="300" swimtime="00:01:33.07" resultid="2387" heatid="4881" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="300" swimtime="00:01:20.69" resultid="2388" heatid="4901" lane="2" entrytime="00:01:19.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="424" swimtime="00:00:30.51" resultid="2389" heatid="5096" lane="6" entrytime="00:00:30.37" entrycourse="SCM" />
                <RESULT eventid="1301" points="299" swimtime="00:00:42.39" resultid="2390" heatid="5042" lane="2" entrytime="00:00:43.49" entrycourse="SCM" />
                <RESULT eventid="4411" points="403" swimtime="00:00:33.00" resultid="5388" heatid="4680" lane="2" />
                <RESULT eventid="4413" points="363" swimtime="00:00:34.16" resultid="5394" heatid="4691" lane="2" />
                <RESULT eventid="5804" points="407" swimtime="00:00:30.94" resultid="10195" heatid="6054" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Kraemer Geremia" birthdate="2011-07-20" gender="F" nation="BRA" license="366908" swrid="5588763" athleteid="2302" externalid="366908" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="326" swimtime="00:00:35.42" resultid="2303" heatid="4657" lane="5" />
                <RESULT eventid="1077" points="404" swimtime="00:00:34.13" resultid="2304" heatid="4722" lane="5" entrytime="00:00:34.61" entrycourse="SCM" />
                <RESULT eventid="1119" points="428" swimtime="00:02:37.80" resultid="2305" heatid="4874" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                    <SPLIT distance="100" swimtime="00:01:58.62" />
                    <SPLIT distance="150" swimtime="00:02:37.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="326" swimtime="00:01:13.00" resultid="2306" heatid="4933" lane="1" entrytime="00:01:06.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="417" swimtime="00:00:30.67" resultid="2307" heatid="5085" lane="2" />
                <RESULT eventid="1301" points="319" swimtime="00:00:41.48" resultid="2308" heatid="5036" lane="8" />
                <RESULT eventid="4411" points="329" swimtime="00:00:35.31" resultid="5356" heatid="4682" lane="4" />
                <RESULT eventid="4413" points="338" swimtime="00:00:34.98" resultid="5361" heatid="4692" lane="3" />
                <RESULT eventid="4417" points="395" swimtime="00:00:34.40" resultid="5426" heatid="4733" lane="1" />
                <RESULT eventid="4419" points="407" swimtime="00:00:34.05" resultid="5433" heatid="4743" lane="1" />
                <RESULT eventid="5801" points="324" swimtime="00:00:41.30" resultid="10160" heatid="6070" lane="6" />
                <RESULT eventid="5804" points="446" swimtime="00:00:30.01" resultid="10200" heatid="6056" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco" lastname="Morais Shibata" birthdate="2014-02-09" gender="M" nation="BRA" license="391018" swrid="5602561" athleteid="2655" externalid="391018" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="82" swimtime="00:00:49.91" resultid="2656" heatid="4754" lane="2" entrytime="00:00:51.40" entrycourse="SCM" />
                <RESULT eventid="1102" points="123" swimtime="00:00:44.34" resultid="2657" heatid="4816" lane="4" entrytime="00:00:43.82" entrycourse="SCM" />
                <RESULT eventid="1213" points="104" swimtime="00:01:57.22" resultid="2658" heatid="4947" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="114" swimtime="00:01:39.66" resultid="2659" heatid="4983" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="103" swimtime="00:00:53.12" resultid="2661" heatid="5128" lane="3" entrytime="00:01:00.68" entrycourse="SCM" />
                <RESULT eventid="4427" points="120" swimtime="00:00:44.75" resultid="5510" heatid="4822" lane="6" />
                <RESULT eventid="10329" points="116" swimtime="00:00:41.26" resultid="10439" heatid="10344" lane="2" entrytime="00:00:39.31" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Baptistella" birthdate="2013-01-23" gender="M" nation="BRA" license="391152" swrid="5602545" athleteid="2725" externalid="391152" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="216" swimtime="00:00:36.24" resultid="2726" heatid="4768" lane="1" />
                <RESULT eventid="1105" points="216" swimtime="00:00:36.85" resultid="2727" heatid="4837" lane="3" entrytime="00:00:38.09" entrycourse="SCM" />
                <RESULT eventid="1249" points="215" swimtime="00:01:20.67" resultid="2728" heatid="4985" lane="2" entrytime="00:01:23.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="243" swimtime="00:01:11.79" resultid="2729" heatid="5003" lane="3" entrytime="00:01:23.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="157" swimtime="00:00:46.21" resultid="2731" heatid="5147" lane="4" />
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente., Na volta dos 25m." eventid="4425" status="DSQ" swimtime="00:00:38.64" resultid="5479" heatid="4804" lane="1" />
                <RESULT eventid="4423" points="218" swimtime="00:00:36.09" resultid="5485" heatid="4792" lane="5" />
                <RESULT eventid="4429" points="218" swimtime="00:00:36.70" resultid="5513" heatid="4852" lane="3" />
                <RESULT eventid="4431" points="207" swimtime="00:00:37.33" resultid="5519" heatid="4864" lane="3" />
                <RESULT eventid="10332" points="263" swimtime="00:00:31.43" resultid="10443" heatid="10349" lane="7" entrytime="00:00:37.09" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Fischer Araujo" birthdate="2013-10-14" gender="M" nation="BRA" license="414420" swrid="5755336" athleteid="3047" externalid="414420" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="24" swimtime="00:01:14.74" resultid="3048" heatid="4771" lane="6" />
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida." eventid="1105" status="DSQ" swimtime="00:00:53.43" resultid="3049" heatid="4830" lane="6" />
                <RESULT eventid="1213" points="66" swimtime="00:02:16.63" resultid="3050" heatid="4948" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="85" swimtime="00:01:41.63" resultid="3051" heatid="4999" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="78" swimtime="00:00:58.38" resultid="3053" heatid="5142" lane="3" />
                <RESULT eventid="10332" points="93" swimtime="00:00:44.38" resultid="10464" heatid="10347" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maya" lastname="Assahida Moreria" birthdate="2014-02-24" gender="F" nation="BRA" license="391020" swrid="5602512" athleteid="2669" externalid="391020" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="143" swimtime="00:00:46.52" resultid="2670" heatid="4651" lane="1" entrytime="00:00:43.73" entrycourse="SCM" />
                <RESULT eventid="1074" points="156" swimtime="00:00:46.90" resultid="2671" heatid="4699" lane="5" entrytime="00:00:54.61" entrycourse="SCM" />
                <RESULT eventid="1165" points="166" swimtime="00:01:39.73" resultid="2672" heatid="4911" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="129" swimtime="00:01:46.72" resultid="2673" heatid="4900" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="167" swimtime="00:00:51.45" resultid="2674" heatid="5025" lane="8" entrytime="00:00:52.64" entrycourse="SCM" />
                <RESULT eventid="1311" points="242" swimtime="00:00:36.77" resultid="2675" heatid="5076" lane="1" entrytime="00:00:38.43" entrycourse="SCM" />
                <RESULT eventid="4439" points="259" swimtime="00:00:35.96" resultid="10184" heatid="6050" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcelo" birthdate="2010-01-09" gender="M" nameprefix="Vanhazebrouck" nation="BRA" license="339043" swrid="5588786" athleteid="10319" externalid="339043" level="CLBO">
              <RESULTS>
                <RESULT eventid="1329" points="326" swimtime="00:00:36.22" resultid="10321" heatid="5137" lane="2" />
                <RESULT eventid="5807" points="330" swimtime="00:00:36.09" resultid="10328" heatid="6042" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Sieczkowski Pacheco" birthdate="2015-11-20" gender="F" nation="BRA" license="393261" swrid="5616450" athleteid="2760" externalid="393261" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="82" swimtime="00:00:55.94" resultid="2761" heatid="4648" lane="5" entrytime="00:01:01.63" entrycourse="SCM" />
                <RESULT eventid="1074" points="96" swimtime="00:00:54.98" resultid="2762" heatid="4700" lane="6" entrytime="00:00:52.41" entrycourse="SCM" />
                <RESULT eventid="1129" points="119" swimtime="00:02:06.69" resultid="2763" heatid="4880" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="94" swimtime="00:02:00.46" resultid="2764" heatid="4908" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="110" swimtime="00:00:59.09" resultid="2765" heatid="5024" lane="1" entrytime="00:00:56.24" entrycourse="SCM" />
                <RESULT eventid="1311" points="153" swimtime="00:00:42.82" resultid="2766" heatid="5072" lane="6" entrytime="00:00:50.99" entrycourse="SCM" />
                <RESULT eventid="4409" points="104" swimtime="00:00:51.74" resultid="5368" heatid="4655" lane="6" />
                <RESULT eventid="4439" points="157" swimtime="00:00:42.50" resultid="10178" heatid="6048" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Jacob Brunetti" birthdate="2015-11-10" gender="M" nation="BRA" license="406837" swrid="5717274" athleteid="2956" externalid="406837" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="29" swimtime="00:01:10.32" resultid="2957" heatid="4752" lane="2" entrytime="00:01:34.76" entrycourse="SCM" />
                <RESULT eventid="1102" points="61" swimtime="00:00:55.98" resultid="2958" heatid="4813" lane="2" entrytime="00:00:59.75" entrycourse="SCM" />
                <RESULT eventid="1213" points="46" swimtime="00:02:33.65" resultid="2959" heatid="4946" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="48" swimtime="00:02:12.76" resultid="2960" heatid="4982" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="48" swimtime="00:01:08.58" resultid="2962" heatid="5127" lane="2" entrytime="00:01:15.32" entrycourse="SCM" />
                <RESULT eventid="10329" points="45" swimtime="00:00:56.49" resultid="10457" heatid="10340" lane="2" entrytime="00:00:59.39" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Taborda Ribas" birthdate="2015-12-30" gender="M" nation="BRA" license="406748" swrid="5717299" athleteid="2921" externalid="406748" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="40" swimtime="00:01:03.39" resultid="2922" heatid="4753" lane="5" entrytime="00:01:26.45" entrycourse="SCM" />
                <RESULT eventid="1102" points="64" swimtime="00:00:55.20" resultid="2923" heatid="4814" lane="6" entrytime="00:00:57.15" entrycourse="SCM" />
                <RESULT eventid="1249" points="68" swimtime="00:01:58.39" resultid="2924" heatid="4981" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="2925" heatid="4997" lane="3" />
                <RESULT eventid="1326" points="52" swimtime="00:01:06.58" resultid="2927" heatid="5127" lane="4" entrytime="00:01:10.29" entrycourse="SCM" />
                <RESULT eventid="10329" points="78" swimtime="00:00:47.16" resultid="10454" heatid="10342" lane="6" entrytime="00:00:48.19" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Zaroni" birthdate="2010-03-03" gender="F" nation="BRA" license="356345" swrid="5600282" athleteid="2197" externalid="356345" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="338" swimtime="00:00:34.98" resultid="2198" heatid="4658" lane="5" />
                <RESULT eventid="1077" points="336" swimtime="00:00:36.32" resultid="2199" heatid="4710" lane="4" />
                <RESULT eventid="1129" points="439" swimtime="00:01:22.02" resultid="2200" heatid="4887" lane="1" entrytime="00:01:22.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="435" swimtime="00:01:06.27" resultid="2201" heatid="4932" lane="4" entrytime="00:01:06.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="360" swimtime="00:00:32.22" resultid="2202" heatid="5094" lane="3" entrytime="00:00:30.88" entrycourse="SCM" />
                <RESULT eventid="1301" points="382" swimtime="00:00:39.09" resultid="2203" heatid="5045" lane="6" entrytime="00:00:38.48" entrycourse="SCM" />
                <RESULT eventid="4411" points="358" swimtime="00:00:34.33" resultid="5328" heatid="4684" lane="3" />
                <RESULT eventid="4413" points="316" swimtime="00:00:35.78" resultid="5334" heatid="4693" lane="3" />
                <RESULT eventid="4417" points="338" swimtime="00:00:36.24" resultid="5436" heatid="4735" lane="1" />
                <RESULT eventid="4419" points="340" swimtime="00:00:36.16" resultid="5442" heatid="4744" lane="1" />
                <RESULT eventid="5801" points="368" swimtime="00:00:39.57" resultid="10105" heatid="6072" lane="3" />
                <RESULT eventid="5804" points="384" swimtime="00:00:31.54" resultid="10209" heatid="6058" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rene" lastname="Osternack Erbe" birthdate="2011-04-03" gender="M" nation="BRA" license="366907" swrid="5588842" athleteid="2295" externalid="366907" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="197" swimtime="00:00:37.36" resultid="2296" heatid="4769" lane="3" />
                <RESULT eventid="1105" points="257" swimtime="00:00:34.77" resultid="2297" heatid="4827" lane="2" />
                <RESULT eventid="1249" points="241" swimtime="00:01:17.60" resultid="2298" heatid="4986" lane="6" entrytime="00:01:18.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1237" points="231" swimtime="00:01:17.80" resultid="2299" heatid="4972" lane="1" entrytime="00:01:29.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="165" swimtime="00:00:45.47" resultid="2301" heatid="5143" lane="5" />
                <RESULT eventid="4429" points="240" swimtime="00:00:35.53" resultid="5575" heatid="4856" lane="6" />
                <RESULT eventid="10332" points="288" swimtime="00:00:30.51" resultid="10410" heatid="10356" lane="7" entrytime="00:00:30.60" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Jarenko Gomes" birthdate="2014-05-17" gender="F" nation="BRA" license="407692" swrid="5725992" athleteid="2997" externalid="407692" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" status="DNS" swimtime="00:00:00.00" resultid="2998" heatid="4647" lane="4" entrytime="00:01:08.17" entrycourse="SCM" />
                <RESULT eventid="1074" status="DNS" swimtime="00:00:00.00" resultid="2999" heatid="4698" lane="6" entrytime="00:00:59.17" entrycourse="SCM" />
                <RESULT eventid="1129" status="DNS" swimtime="00:00:00.00" resultid="3000" heatid="4882" lane="4" />
                <RESULT eventid="1189" status="DNS" swimtime="00:00:00.00" resultid="3001" heatid="4924" lane="4" />
                <RESULT eventid="1298" status="DNS" swimtime="00:00:00.00" resultid="3002" heatid="5023" lane="1" entrytime="00:01:02.82" entrycourse="SCM" />
                <RESULT eventid="1311" status="DNS" swimtime="00:00:00.00" resultid="3003" heatid="5071" lane="2" entrytime="00:00:52.18" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Clara Prado Biscaia" birthdate="2013-10-24" gender="F" nation="BRA" license="391015" swrid="5602526" athleteid="2643" externalid="391015" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="194" swimtime="00:00:42.10" resultid="2644" heatid="4667" lane="2" entrytime="00:00:43.81" entrycourse="SCM" />
                <RESULT eventid="1077" points="157" swimtime="00:00:46.77" resultid="2645" heatid="4715" lane="6" entrytime="00:00:51.80" entrycourse="SCM" />
                <RESULT eventid="1314" points="248" swimtime="00:00:36.49" resultid="2646" heatid="5088" lane="8" entrytime="00:00:37.59" entrycourse="SCM" />
                <RESULT eventid="1301" points="134" swimtime="00:00:55.31" resultid="2647" heatid="5040" lane="7" entrytime="00:00:58.39" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Cabrera Cirino" birthdate="2011-01-28" gender="M" nation="BRA" license="369531" swrid="5588569" athleteid="2419" externalid="369531" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="372" swimtime="00:00:30.23" resultid="2420" heatid="4774" lane="6" />
                <RESULT eventid="1105" points="349" swimtime="00:00:31.38" resultid="2421" heatid="4833" lane="5" />
                <RESULT eventid="1227" points="451" swimtime="00:02:09.55" resultid="2422" heatid="4964" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                    <SPLIT distance="100" swimtime="00:01:03.10" />
                    <SPLIT distance="150" swimtime="00:01:36.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="428" swimtime="00:00:59.50" resultid="2423" heatid="5009" lane="6" entrytime="00:01:01.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" status="DNS" swimtime="00:00:00.00" resultid="2425" heatid="5138" lane="5" />
                <RESULT eventid="4423" points="361" swimtime="00:00:30.53" resultid="5530" heatid="4796" lane="2" />
                <RESULT eventid="4425" points="298" swimtime="00:00:32.53" resultid="5536" heatid="4806" lane="2" />
                <RESULT eventid="4429" points="344" swimtime="00:00:31.53" resultid="5566" heatid="4856" lane="1" />
                <RESULT eventid="4431" points="340" swimtime="00:00:31.65" resultid="5572" heatid="4866" lane="1" />
                <RESULT eventid="10332" points="424" swimtime="00:00:26.82" resultid="10421" heatid="10357" lane="4" entrytime="00:00:28.24" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Lazzarotti Matias" birthdate="2012-03-19" gender="F" nation="BRA" license="391026" swrid="5602552" athleteid="2704" externalid="391026" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="284" swimtime="00:00:37.05" resultid="2705" heatid="4657" lane="2" />
                <RESULT eventid="1077" points="372" swimtime="00:00:35.10" resultid="2706" heatid="4722" lane="1" entrytime="00:00:34.84" entrycourse="SCM" />
                <RESULT eventid="1165" points="348" swimtime="00:01:17.99" resultid="2707" heatid="4914" lane="6" entrytime="00:01:17.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="388" swimtime="00:02:31.21" resultid="2708" heatid="4894" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                    <SPLIT distance="100" swimtime="00:01:15.58" />
                    <SPLIT distance="150" swimtime="00:01:54.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="375" swimtime="00:00:31.77" resultid="2709" heatid="5093" lane="8" entrytime="00:00:32.63" entrycourse="SCM" />
                <RESULT eventid="1301" points="272" swimtime="00:00:43.74" resultid="2710" heatid="5044" lane="7" entrytime="00:00:42.49" entrycourse="SCM" />
                <RESULT eventid="4417" points="333" swimtime="00:00:36.41" resultid="5419" heatid="4731" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Carneiro Silva" birthdate="2011-02-21" gender="F" nation="BRA" license="390924" swrid="5602522" athleteid="2865" externalid="390924" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="301" swimtime="00:00:36.35" resultid="2866" heatid="4664" lane="4" />
                <RESULT eventid="1077" points="317" swimtime="00:00:37.03" resultid="2867" heatid="4721" lane="6" entrytime="00:00:36.94" entrycourse="SCM" />
                <RESULT eventid="1143" points="367" swimtime="00:02:34.00" resultid="2868" heatid="4893" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="359" swimtime="00:01:10.66" resultid="2869" heatid="4931" lane="5" entrytime="00:01:11.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="378" swimtime="00:00:31.70" resultid="2870" heatid="5092" lane="5" entrytime="00:00:32.92" entrycourse="SCM" />
                <RESULT eventid="1301" points="279" swimtime="00:00:43.37" resultid="2871" heatid="5036" lane="5" />
                <RESULT eventid="5804" points="361" swimtime="00:00:32.20" resultid="10203" heatid="6056" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Coelho" birthdate="2011-11-11" gender="M" nation="BRA" license="366889" swrid="5602527" athleteid="2239" externalid="366889" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="307" swimtime="00:00:32.23" resultid="2240" heatid="4769" lane="6" />
                <RESULT eventid="1105" points="201" swimtime="00:00:37.71" resultid="2241" heatid="4826" lane="5" />
                <RESULT comment="SW 7.5 - Executou uma pernada de borboleta durante o nado.  (Horário: 1:03)" eventid="1213" status="DSQ" swimtime="00:01:25.48" resultid="2242" heatid="4951" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1237" points="251" swimtime="00:01:15.71" resultid="2243" heatid="4973" lane="4" entrytime="00:01:14.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="252" swimtime="00:00:39.49" resultid="2245" heatid="5142" lane="5" />
                <RESULT eventid="4423" points="285" swimtime="00:00:33.05" resultid="5534" heatid="4796" lane="6" />
                <RESULT eventid="10332" points="304" swimtime="00:00:29.98" resultid="10406" heatid="10348" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Portes Fabiane" birthdate="2012-12-28" gender="M" nation="BRA" license="376983" swrid="5588864" athleteid="2503" externalid="376983" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="63" swimtime="00:00:54.45" resultid="2504" heatid="4763" lane="3" />
                <RESULT eventid="1105" points="74" swimtime="00:00:52.62" resultid="2505" heatid="4834" lane="4" entrytime="00:00:51.36" entrycourse="SCM" />
                <RESULT eventid="1249" points="81" swimtime="00:01:51.46" resultid="2506" heatid="4984" lane="6" entrytime="00:01:52.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="111" swimtime="00:01:33.26" resultid="2507" heatid="5002" lane="5" entrytime="00:01:38.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="88" swimtime="00:00:55.90" resultid="2509" heatid="5148" lane="2" entrytime="00:00:59.61" entrycourse="SCM" />
                <RESULT eventid="10332" points="111" swimtime="00:00:41.85" resultid="10425" heatid="10349" lane="1" entrytime="00:00:45.07" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luigi" lastname="Antoniuk Paganini" birthdate="2014-11-13" gender="M" nation="BRA" license="382127" swrid="5602509" athleteid="2587" externalid="382127" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="130" swimtime="00:00:42.88" resultid="2588" heatid="4756" lane="6" entrytime="00:00:43.75" entrycourse="SCM" />
                <RESULT eventid="1102" points="146" swimtime="00:00:41.94" resultid="2589" heatid="4817" lane="1" entrytime="00:00:42.68" entrycourse="SCM" />
                <RESULT eventid="1249" points="140" swimtime="00:01:32.86" resultid="2590" heatid="4981" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1237" points="123" swimtime="00:01:35.98" resultid="2591" heatid="4971" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="95" swimtime="00:00:54.49" resultid="2593" heatid="5131" lane="7" entrytime="00:00:54.89" entrycourse="SCM" />
                <RESULT eventid="4421" points="133" swimtime="00:00:42.53" resultid="5474" heatid="4761" lane="6" />
                <RESULT eventid="4427" points="148" swimtime="00:00:41.76" resultid="5508" heatid="4822" lane="4" />
                <RESULT eventid="10329" points="184" swimtime="00:00:35.40" resultid="10433" heatid="10345" lane="6" entrytime="00:00:36.20" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Prosdocimo" birthdate="2012-11-30" gender="M" nation="BRA" license="369272" swrid="5602575" athleteid="2363" externalid="369272" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="213" swimtime="00:00:36.40" resultid="2364" heatid="4776" lane="4" entrytime="00:00:38.13" entrycourse="SCM" />
                <RESULT eventid="1105" points="220" swimtime="00:00:36.59" resultid="2365" heatid="4838" lane="2" entrytime="00:00:37.07" entrycourse="SCM" />
                <RESULT eventid="1203" points="257" swimtime="00:02:46.06" resultid="2366" heatid="4942" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.62" />
                    <SPLIT distance="100" swimtime="00:01:21.08" />
                    <SPLIT distance="150" swimtime="00:02:03.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="283" swimtime="00:01:08.25" resultid="2367" heatid="5007" lane="2" entrytime="00:01:07.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="149" swimtime="00:00:47.05" resultid="2369" heatid="5146" lane="8" />
                <RESULT eventid="4429" points="225" swimtime="00:00:36.33" resultid="5524" heatid="4854" lane="5" />
                <RESULT eventid="10332" points="274" swimtime="00:00:31.02" resultid="10417" heatid="10355" lane="4" entrytime="00:00:30.90" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Cavalca Petraglia" birthdate="2015-08-06" gender="M" nation="BRA" license="397275" swrid="5641757" athleteid="2816" externalid="397275" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="78" swimtime="00:00:50.77" resultid="2817" heatid="4754" lane="4" entrytime="00:00:51.02" entrycourse="SCM" />
                <RESULT eventid="1102" points="80" swimtime="00:00:51.31" resultid="2818" heatid="4815" lane="5" entrytime="00:00:50.39" entrycourse="SCM" />
                <RESULT eventid="1213" points="85" swimtime="00:02:05.60" resultid="2819" heatid="4950" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1237" points="55" swimtime="00:02:05.29" resultid="2820" heatid="4969" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="82" swimtime="00:00:57.23" resultid="2822" heatid="5130" lane="1" entrytime="00:00:58.05" entrycourse="SCM" />
                <RESULT eventid="10329" points="91" swimtime="00:00:44.69" resultid="10448" heatid="10342" lane="2" entrytime="00:00:44.65" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorena" lastname="Mascarenhas" birthdate="2011-08-31" gender="F" nation="BRA" license="370581" swrid="5602558" athleteid="2447" externalid="370581" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="319" swimtime="00:00:35.66" resultid="2448" heatid="4666" lane="6" />
                <RESULT eventid="1077" points="363" swimtime="00:00:35.39" resultid="2449" heatid="4721" lane="2" entrytime="00:00:35.97" entrycourse="SCM" />
                <RESULT eventid="1165" points="412" swimtime="00:01:13.75" resultid="2450" heatid="4914" lane="5" entrytime="00:01:16.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="383" swimtime="00:01:09.14" resultid="2451" heatid="4931" lane="1" entrytime="00:01:11.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="395" swimtime="00:00:31.23" resultid="2452" heatid="5083" lane="3" />
                <RESULT eventid="1301" points="384" swimtime="00:00:39.01" resultid="2453" heatid="5044" lane="2" entrytime="00:00:40.17" entrycourse="SCM" />
                <RESULT eventid="4411" points="314" swimtime="00:00:35.85" resultid="5358" heatid="4682" lane="6" />
                <RESULT eventid="4417" points="375" swimtime="00:00:34.99" resultid="5432" heatid="4733" lane="2" />
                <RESULT eventid="4419" points="370" swimtime="00:00:35.17" resultid="5434" heatid="4743" lane="2" />
                <RESULT eventid="5801" points="358" swimtime="00:00:39.94" resultid="10156" heatid="6070" lane="3" />
                <RESULT eventid="5804" points="408" swimtime="00:00:30.90" resultid="10199" heatid="6056" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joana" lastname="Asinelli Casagrande" birthdate="2013-10-26" gender="F" nation="BRA" license="376970" swrid="5588536" athleteid="2482" externalid="376970" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="262" swimtime="00:00:38.06" resultid="2483" heatid="4668" lane="4" entrytime="00:00:39.22" entrycourse="SCM" />
                <RESULT eventid="1077" points="305" swimtime="00:00:37.49" resultid="2484" heatid="4719" lane="2" entrytime="00:00:39.31" entrycourse="SCM" />
                <RESULT eventid="1119" points="301" swimtime="00:02:57.38" resultid="2485" heatid="4874" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.95" />
                    <SPLIT distance="100" swimtime="00:02:12.60" />
                    <SPLIT distance="150" swimtime="00:02:57.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="305" swimtime="00:01:21.53" resultid="2486" heatid="4913" lane="1" entrytime="00:01:24.94" entrycourse="SCM" />
                <RESULT eventid="1314" points="315" swimtime="00:00:33.70" resultid="2487" heatid="5086" lane="2" entrytime="00:00:39.14" entrycourse="SCM" />
                <RESULT eventid="1301" points="209" swimtime="00:00:47.77" resultid="2488" heatid="5041" lane="8" entrytime="00:00:53.15" entrycourse="SCM" />
                <RESULT eventid="4417" points="307" swimtime="00:00:37.41" resultid="5408" heatid="4729" lane="1" />
                <RESULT eventid="4419" points="285" swimtime="00:00:38.36" resultid="5414" heatid="4741" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Betina" lastname="Vieira Pellanda" birthdate="2014-02-16" gender="F" nation="BRA" license="391041" swrid="5602589" athleteid="2718" externalid="391041" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="137" swimtime="00:00:47.25" resultid="2719" heatid="4648" lane="1" entrytime="00:01:01.99" entrycourse="SCM" />
                <RESULT eventid="1074" points="151" swimtime="00:00:47.41" resultid="2720" heatid="4701" lane="1" entrytime="00:00:49.00" entrycourse="SCM" />
                <RESULT eventid="1129" points="176" swimtime="00:01:51.21" resultid="2721" heatid="4879" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="127" swimtime="00:01:48.98" resultid="2722" heatid="4906" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="168" swimtime="00:00:51.41" resultid="2723" heatid="5024" lane="6" entrytime="00:00:56.10" entrycourse="SCM" />
                <RESULT eventid="1311" points="195" swimtime="00:00:39.50" resultid="2724" heatid="5073" lane="8" entrytime="00:00:42.42" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ravi" lastname="Osternack Erbe" birthdate="2013-08-10" gender="M" nation="BRA" license="372681" swrid="5588841" athleteid="2426" externalid="372681" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="205" swimtime="00:00:36.83" resultid="2427" heatid="4778" lane="6" entrytime="00:00:35.96" entrycourse="SCM" />
                <RESULT eventid="1105" points="139" swimtime="00:00:42.66" resultid="2428" heatid="4836" lane="2" entrytime="00:00:40.46" entrycourse="SCM" />
                <RESULT eventid="1237" points="177" swimtime="00:01:25.09" resultid="2429" heatid="4972" lane="4" entrytime="00:01:24.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="203" swimtime="00:01:16.24" resultid="2430" heatid="5006" lane="2" entrytime="00:01:12.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.1 - Mais de uma pernada de borboleta antes da primeira pernada de peito após o início ou a virada., Após a  volta dos 25m." eventid="1329" status="DSQ" swimtime="00:00:43.06" resultid="2432" heatid="5151" lane="8" entrytime="00:00:47.13" entrycourse="SCM" />
                <RESULT eventid="4423" points="217" swimtime="00:00:36.18" resultid="5486" heatid="4792" lane="6" />
                <RESULT eventid="10332" points="200" swimtime="00:00:34.44" resultid="10422" heatid="10353" lane="2" entrytime="00:00:32.82" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Antunes Luzzi" birthdate="2014-02-14" gender="M" nation="BRA" license="391019" swrid="5602510" athleteid="2662" externalid="391019" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="33" swimtime="00:01:07.64" resultid="2663" heatid="4752" lane="4" entrytime="00:01:34.31" entrycourse="SCM" />
                <RESULT eventid="1102" points="44" swimtime="00:01:02.26" resultid="2664" heatid="4813" lane="3" entrytime="00:00:57.61" entrycourse="SCM" />
                <RESULT eventid="1249" points="60" swimtime="00:02:02.82" resultid="2665" heatid="4981" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="57" swimtime="00:01:56.49" resultid="2666" heatid="4996" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="68" swimtime="00:01:00.98" resultid="2668" heatid="5130" lane="7" entrytime="00:00:59.82" entrycourse="SCM" />
                <RESULT eventid="10329" status="DNS" swimtime="00:00:00.00" resultid="10440" heatid="10342" lane="7" entrytime="00:00:49.66" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Cipriani Presiazniuk" birthdate="2012-07-03" gender="M" nation="BRA" license="369267" swrid="5588594" athleteid="2337" externalid="369267" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="188" swimtime="00:00:37.93" resultid="2338" heatid="4771" lane="3" />
                <RESULT eventid="1105" points="207" swimtime="00:00:37.36" resultid="2339" heatid="4838" lane="5" entrytime="00:00:37.28" entrycourse="SCM" />
                <RESULT eventid="1203" points="226" swimtime="00:02:53.37" resultid="2340" heatid="4943" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.93" />
                    <SPLIT distance="100" swimtime="00:01:27.64" />
                    <SPLIT distance="150" swimtime="00:02:12.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="209" swimtime="00:01:21.39" resultid="2341" heatid="4985" lane="3" entrytime="00:01:22.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="171" swimtime="00:00:44.92" resultid="2343" heatid="5143" lane="3" />
                <RESULT eventid="4429" points="210" swimtime="00:00:37.15" resultid="5525" heatid="4854" lane="6" />
                <RESULT eventid="10332" points="271" swimtime="00:00:31.12" resultid="10413" heatid="10352" lane="8" entrytime="00:00:32.90" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="De Fortes" birthdate="2015-06-01" gender="M" nation="BRA" license="399680" swrid="5652884" athleteid="2830" externalid="399680" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="100" swimtime="00:00:46.80" resultid="2831" heatid="4755" lane="5" entrytime="00:00:46.93" entrycourse="SCM" />
                <RESULT eventid="1102" points="97" swimtime="00:00:47.99" resultid="2832" heatid="4816" lane="1" entrytime="00:00:48.02" entrycourse="SCM" />
                <RESULT eventid="1249" status="DNS" swimtime="00:00:00.00" resultid="2833" heatid="4981" lane="5" />
                <RESULT eventid="1237" status="DNS" swimtime="00:00:00.00" resultid="2834" heatid="4970" lane="6" />
                <RESULT eventid="1326" status="DNS" swimtime="00:00:00.00" resultid="2836" heatid="5126" lane="6" />
                <RESULT eventid="4421" points="115" swimtime="00:00:44.71" resultid="5467" heatid="4760" lane="5" />
                <RESULT eventid="10329" status="DNS" swimtime="00:00:00.00" resultid="10449" heatid="10344" lane="6" entrytime="00:00:38.66" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Vian" birthdate="2014-03-25" gender="F" nation="BRA" license="393919" swrid="5641779" athleteid="2795" externalid="393919" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="134" swimtime="00:00:47.56" resultid="2796" heatid="4650" lane="2" entrytime="00:00:48.99" entrycourse="SCM" />
                <RESULT eventid="1074" points="187" swimtime="00:00:44.14" resultid="2797" heatid="4702" lane="6" entrytime="00:00:47.99" entrycourse="SCM" />
                <RESULT eventid="1165" points="157" swimtime="00:01:41.62" resultid="2798" heatid="4908" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="163" swimtime="00:01:31.89" resultid="2799" heatid="4927" lane="6" entrytime="00:01:42.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="101" swimtime="00:01:00.89" resultid="2800" heatid="5023" lane="4" entrytime="00:00:59.76" entrycourse="SCM" />
                <RESULT eventid="1311" points="190" swimtime="00:00:39.87" resultid="2801" heatid="5073" lane="7" entrytime="00:00:42.69" entrycourse="SCM" />
                <RESULT eventid="4415" points="186" swimtime="00:00:44.22" resultid="5405" heatid="4707" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolau" lastname="Neto" birthdate="2011-03-22" gender="M" nation="BRA" license="366906" swrid="5602565" athleteid="2288" externalid="366906" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="224" swimtime="00:00:35.79" resultid="2289" heatid="4774" lane="4" />
                <RESULT eventid="1105" points="178" swimtime="00:00:39.30" resultid="2290" heatid="4833" lane="6" />
                <RESULT eventid="1213" points="386" swimtime="00:01:15.89" resultid="2291" heatid="4953" lane="4" entrytime="00:01:22.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="330" swimtime="00:02:53.79" resultid="2292" heatid="4993" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                    <SPLIT distance="100" swimtime="00:01:24.21" />
                    <SPLIT distance="150" swimtime="00:02:08.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="345" swimtime="00:00:35.54" resultid="2294" heatid="5152" lane="3" entrytime="00:00:40.50" entrycourse="SCM" />
                <RESULT eventid="5807" points="359" swimtime="00:00:35.10" resultid="10282" heatid="6040" lane="5" />
                <RESULT eventid="10332" points="358" swimtime="00:00:28.37" resultid="10409" heatid="10357" lane="8" entrytime="00:00:29.70" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Albuquerque" birthdate="2012-11-16" gender="F" nation="BRA" license="369281" swrid="5602506" athleteid="2405" externalid="369281" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="268" swimtime="00:00:37.79" resultid="2406" heatid="4669" lane="2" entrytime="00:00:38.36" entrycourse="SCM" />
                <RESULT eventid="1077" points="281" swimtime="00:00:38.53" resultid="2407" heatid="4718" lane="1" entrytime="00:00:41.18" entrycourse="SCM" />
                <RESULT eventid="1129" points="345" swimtime="00:01:28.84" resultid="2408" heatid="4886" lane="5" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="350" swimtime="00:03:10.80" resultid="2409" heatid="4921" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.44" />
                    <SPLIT distance="100" swimtime="00:01:33.85" />
                    <SPLIT distance="150" swimtime="00:02:22.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="336" swimtime="00:00:32.98" resultid="2410" heatid="5084" lane="6" />
                <RESULT eventid="1301" points="333" swimtime="00:00:40.89" resultid="2411" heatid="5045" lane="8" entrytime="00:00:41.79" entrycourse="SCM" />
                <RESULT eventid="5801" points="333" swimtime="00:00:40.90" resultid="10101" heatid="6068" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Pereira Galle" birthdate="2011-08-02" gender="F" nation="BRA" license="369465" swrid="5627330" athleteid="2872" externalid="369465" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="326" swimtime="00:00:35.39" resultid="2873" heatid="4663" lane="1" />
                <RESULT eventid="1077" points="243" swimtime="00:00:40.46" resultid="2874" heatid="4708" lane="3" />
                <RESULT eventid="1129" points="365" swimtime="00:01:27.24" resultid="2875" heatid="4886" lane="2" entrytime="00:01:26.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="370" swimtime="00:01:09.96" resultid="2876" heatid="4932" lane="1" entrytime="00:01:08.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="365" swimtime="00:00:32.06" resultid="2877" heatid="5084" lane="5" />
                <RESULT eventid="1301" points="396" swimtime="00:00:38.62" resultid="2878" heatid="5038" lane="2" />
                <RESULT eventid="4411" points="320" swimtime="00:00:35.61" resultid="5355" heatid="4682" lane="3" />
                <RESULT eventid="5801" points="414" swimtime="00:00:38.04" resultid="10155" heatid="6070" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gael" lastname="Stramandinoli Zanicotti" birthdate="2015-03-21" gender="M" nation="BRA" license="406954" swrid="5717298" athleteid="2970" externalid="406954" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" status="DNS" swimtime="00:00:00.00" resultid="2971" heatid="4753" lane="6" entrytime="00:01:31.38" entrycourse="SCM" />
                <RESULT eventid="1102" status="DNS" swimtime="00:00:00.00" resultid="2972" heatid="4813" lane="6" entrytime="00:01:03.19" entrycourse="SCM" />
                <RESULT eventid="1249" status="DNS" swimtime="00:00:00.00" resultid="2973" heatid="4978" lane="5" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="2974" heatid="5001" lane="5" entrytime="00:02:10.99" entrycourse="SCM" />
                <RESULT eventid="1326" status="DNS" swimtime="00:00:00.00" resultid="2976" heatid="5126" lane="3" entrytime="00:01:32.93" entrycourse="SCM" />
                <RESULT eventid="10329" status="DNS" swimtime="00:00:00.00" resultid="10458" heatid="10341" lane="4" entrytime="00:00:54.87" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Emili Gomes Xavier" birthdate="2010-09-08" gender="F" nation="BRA" license="372519" swrid="5717260" athleteid="2190" externalid="372519" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="322" swimtime="00:00:35.55" resultid="2191" heatid="4662" lane="4" />
                <RESULT eventid="1077" points="323" swimtime="00:00:36.79" resultid="2192" heatid="4721" lane="5" entrytime="00:00:36.12" entrycourse="SCM" />
                <RESULT eventid="1119" points="356" swimtime="00:02:47.74" resultid="2193" heatid="4874" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                    <SPLIT distance="100" swimtime="00:02:05.95" />
                    <SPLIT distance="150" swimtime="00:02:47.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="287" swimtime="00:01:21.94" resultid="2194" heatid="4900" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="451" swimtime="00:00:29.90" resultid="2195" heatid="5085" lane="6" />
                <RESULT eventid="1301" points="414" swimtime="00:00:38.05" resultid="2196" heatid="5045" lane="1" entrytime="00:00:38.19" entrycourse="SCM" />
                <RESULT eventid="4411" points="330" swimtime="00:00:35.27" resultid="5329" heatid="4684" lane="4" />
                <RESULT eventid="4417" points="334" swimtime="00:00:36.37" resultid="5438" heatid="4735" lane="3" />
                <RESULT eventid="4419" points="317" swimtime="00:00:37.00" resultid="5444" heatid="4744" lane="3" />
                <RESULT eventid="5801" points="381" swimtime="00:00:39.10" resultid="10108" heatid="6072" lane="6" />
                <RESULT eventid="5804" points="468" swimtime="00:00:29.52" resultid="10207" heatid="6058" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giulia" lastname="Ziliotto Mehl" birthdate="2015-10-09" gender="F" nation="BRA" license="400122" swrid="5652905" athleteid="2851" externalid="400122" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" status="DNS" swimtime="00:00:00.00" resultid="2852" heatid="4648" lane="3" entrytime="00:00:56.49" entrycourse="SCM" />
                <RESULT eventid="1074" status="DNS" swimtime="00:00:00.00" resultid="2853" heatid="4696" lane="2" />
                <RESULT eventid="1129" status="DNS" swimtime="00:00:00.00" resultid="2854" heatid="4880" lane="3" />
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="2855" heatid="4907" lane="4" />
                <RESULT eventid="1298" status="DNS" swimtime="00:00:00.00" resultid="2856" heatid="5024" lane="5" entrytime="00:00:56.00" entrycourse="SCM" />
                <RESULT eventid="1311" status="DNS" swimtime="00:00:00.00" resultid="2857" heatid="5075" lane="5" entrytime="00:00:42.02" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Rossi Mattioli" birthdate="2013-05-08" gender="F" nation="BRA" license="376988" swrid="5588892" athleteid="2545" externalid="376988" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="259" swimtime="00:00:38.20" resultid="2546" heatid="4665" lane="3" />
                <RESULT eventid="1077" points="290" swimtime="00:00:38.12" resultid="2547" heatid="4719" lane="4" entrytime="00:00:39.12" entrycourse="SCM" />
                <RESULT eventid="1129" points="279" swimtime="00:01:35.42" resultid="2548" heatid="4885" lane="5" entrytime="00:01:39.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="252" swimtime="00:03:33.03" resultid="2549" heatid="4921" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.93" />
                    <SPLIT distance="100" swimtime="00:01:40.88" />
                    <SPLIT distance="150" swimtime="00:02:37.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="315" swimtime="00:00:33.68" resultid="2550" heatid="5092" lane="8" entrytime="00:00:33.29" entrycourse="SCM" />
                <RESULT eventid="1301" points="325" swimtime="00:00:41.23" resultid="2551" heatid="5041" lane="5" entrytime="00:00:47.29" entrycourse="SCM" />
                <RESULT eventid="4417" points="319" swimtime="00:00:36.93" resultid="5409" heatid="4729" lane="2" />
                <RESULT eventid="4419" points="269" swimtime="00:00:39.10" resultid="5415" heatid="4741" lane="2" />
                <RESULT eventid="5801" points="326" swimtime="00:00:41.21" resultid="10092" heatid="6066" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Almeida Jorge" birthdate="2015-05-27" gender="M" nation="BRA" license="406836" swrid="5717242" athleteid="2949" externalid="406836" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="39" swimtime="00:01:03.84" resultid="2950" heatid="4753" lane="2" entrytime="00:01:17.22" entrycourse="SCM" />
                <RESULT eventid="1102" points="65" swimtime="00:00:54.85" resultid="2951" heatid="4810" lane="4" />
                <RESULT eventid="1213" points="82" swimtime="00:02:07.14" resultid="2952" heatid="4950" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="59" swimtime="00:02:03.67" resultid="2953" heatid="4980" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="88" swimtime="00:00:55.93" resultid="2955" heatid="5128" lane="1" entrytime="00:01:02.96" entrycourse="SCM" />
                <RESULT eventid="4445" points="93" swimtime="00:00:55.04" resultid="10311" heatid="6032" lane="7" />
                <RESULT eventid="10329" points="51" swimtime="00:00:54.05" resultid="10456" heatid="10340" lane="4" entrytime="00:00:58.30" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cecilia" lastname="Cabrini Vieira" birthdate="2012-02-11" gender="F" nation="BRA" license="376961" swrid="5588571" athleteid="2468" externalid="376961" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="294" swimtime="00:00:36.65" resultid="2469" heatid="4670" lane="6" entrytime="00:00:38.10" entrycourse="SCM" />
                <RESULT eventid="1077" points="360" swimtime="00:00:35.49" resultid="2470" heatid="4722" lane="6" entrytime="00:00:35.14" entrycourse="SCM" />
                <RESULT eventid="1143" points="442" swimtime="00:02:24.77" resultid="2471" heatid="4895" lane="4" entrytime="00:02:31.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                    <SPLIT distance="100" swimtime="00:01:10.42" />
                    <SPLIT distance="150" swimtime="00:01:48.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="434" swimtime="00:01:06.32" resultid="2472" heatid="4933" lane="6" entrytime="00:01:06.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="423" swimtime="00:00:30.54" resultid="2473" heatid="5097" lane="8" entrytime="00:00:30.03" entrycourse="SCM" />
                <RESULT eventid="1301" points="251" swimtime="00:00:44.93" resultid="2474" heatid="5037" lane="3" />
                <RESULT eventid="4417" points="307" swimtime="00:00:37.40" resultid="5420" heatid="4731" lane="4" />
                <RESULT eventid="5804" points="424" swimtime="00:00:30.52" resultid="10193" heatid="6054" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Livia Bittencourt" birthdate="2015-11-23" gender="F" nation="BRA" license="393260" swrid="5616446" athleteid="2753" externalid="393260" level="CLBO">
              <RESULTS>
                <RESULT comment="SW 8.3 - Movimento de pernada de peito.&#10;&#10;&#10;&#10;&#10;&#10;&#10;" eventid="1061" status="DSQ" swimtime="00:01:04.46" resultid="2754" heatid="4647" lane="2" entrytime="00:01:11.43" entrycourse="SCM" />
                <RESULT eventid="1074" points="78" swimtime="00:00:58.90" resultid="2755" heatid="4698" lane="5" entrytime="00:00:57.18" entrycourse="SCM" />
                <RESULT eventid="1129" points="106" swimtime="00:02:11.54" resultid="2756" heatid="4880" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="2757" heatid="4905" lane="2" />
                <RESULT eventid="1298" points="103" swimtime="00:01:00.50" resultid="2758" heatid="5023" lane="8" entrytime="00:01:03.47" entrycourse="SCM" />
                <RESULT eventid="1311" points="85" swimtime="00:00:52.14" resultid="2759" heatid="5071" lane="7" entrytime="00:01:01.13" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Massimo" lastname="Puppi Cardoso" birthdate="2015-03-30" gender="M" nation="BRA" license="406742" swrid="5717290" athleteid="2893" externalid="406742" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" status="DNS" swimtime="00:00:00.00" resultid="2894" heatid="4753" lane="4" entrytime="00:01:13.69" entrycourse="SCM" />
                <RESULT eventid="1102" status="DNS" swimtime="00:00:00.00" resultid="2895" heatid="4814" lane="1" entrytime="00:00:56.98" entrycourse="SCM" />
                <RESULT eventid="1213" status="DNS" swimtime="00:00:00.00" resultid="2896" heatid="4951" lane="5" />
                <RESULT eventid="1249" status="DNS" swimtime="00:00:00.00" resultid="2897" heatid="4982" lane="1" />
                <RESULT eventid="1326" status="DNS" swimtime="00:00:00.00" resultid="2899" heatid="5130" lane="2" entrytime="00:00:58.72" entrycourse="SCM" />
                <RESULT eventid="10329" status="DNS" swimtime="00:00:00.00" resultid="10452" heatid="10341" lane="6" entrytime="00:00:55.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Leal Souza" birthdate="2014-12-30" gender="M" nation="BRA" license="420717" athleteid="3072" externalid="420717" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="39" swimtime="00:01:03.67" resultid="3073" heatid="4752" lane="6" />
                <RESULT eventid="1102" points="55" swimtime="00:00:57.89" resultid="3074" heatid="4811" lane="5" />
                <RESULT eventid="1213" points="54" swimtime="00:02:25.50" resultid="3075" heatid="4948" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="57" swimtime="00:01:56.13" resultid="3076" heatid="4996" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="47" swimtime="00:01:08.99" resultid="3078" heatid="5126" lane="7" />
                <RESULT eventid="10329" points="70" swimtime="00:00:48.77" resultid="10468" heatid="10341" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Petraglia" birthdate="2012-03-28" gender="M" nation="BRA" license="369282" swrid="5602569" athleteid="2412" externalid="369282" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="146" swimtime="00:00:41.28" resultid="2413" heatid="4771" lane="5" />
                <RESULT eventid="1105" points="183" swimtime="00:00:38.90" resultid="2414" heatid="4837" lane="5" entrytime="00:00:38.74" entrycourse="SCM" />
                <RESULT eventid="1203" points="208" swimtime="00:02:58.03" resultid="2415" heatid="4943" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.16" />
                    <SPLIT distance="100" swimtime="00:01:28.35" />
                    <SPLIT distance="150" swimtime="00:02:14.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="255" swimtime="00:01:10.64" resultid="2416" heatid="5005" lane="1" entrytime="00:01:16.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="193" swimtime="00:00:43.15" resultid="2418" heatid="5152" lane="5" entrytime="00:00:42.44" entrycourse="SCM" />
                <RESULT eventid="10332" points="238" swimtime="00:00:32.49" resultid="10420" heatid="10353" lane="7" entrytime="00:00:33.30" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nina" lastname="Rocha Ribeiro Da Silva" birthdate="2010-09-22" gender="F" nation="BRA" license="367216" swrid="5588884" athleteid="2601" externalid="367216" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="356" swimtime="00:00:34.37" resultid="2602" heatid="4658" lane="4" />
                <RESULT eventid="1077" points="264" swimtime="00:00:39.33" resultid="2603" heatid="4711" lane="5" />
                <RESULT eventid="1129" points="479" swimtime="00:01:19.65" resultid="2604" heatid="4887" lane="4" entrytime="00:01:20.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="422" swimtime="00:01:06.96" resultid="2605" heatid="4932" lane="2" entrytime="00:01:07.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="429" swimtime="00:00:30.38" resultid="2606" heatid="5096" lane="8" entrytime="00:00:30.76" entrycourse="SCM" />
                <RESULT eventid="1301" points="478" swimtime="00:00:36.27" resultid="2607" heatid="5045" lane="4" entrytime="00:00:36.67" entrycourse="SCM" />
                <RESULT eventid="4411" points="358" swimtime="00:00:34.31" resultid="5326" heatid="4684" lane="1" />
                <RESULT eventid="4413" points="303" swimtime="00:00:36.27" resultid="5332" heatid="4693" lane="1" />
                <RESULT eventid="4417" points="264" swimtime="00:00:39.32" resultid="5441" heatid="4735" lane="6" />
                <RESULT eventid="5801" points="480" swimtime="00:00:36.23" resultid="10103" heatid="6072" lane="1" />
                <RESULT eventid="5804" points="440" swimtime="00:00:30.14" resultid="10205" heatid="6058" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Moreira Pasqual" birthdate="2014-07-09" gender="M" nation="BRA" license="382125" swrid="5602562" athleteid="2580" externalid="382125" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="143" swimtime="00:00:41.57" resultid="2581" heatid="4756" lane="5" entrytime="00:00:41.87" entrycourse="SCM" />
                <RESULT eventid="1102" points="114" swimtime="00:00:45.53" resultid="2582" heatid="4816" lane="5" entrytime="00:00:46.42" entrycourse="SCM" />
                <RESULT eventid="1213" points="143" swimtime="00:01:45.51" resultid="2583" heatid="4949" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="107" swimtime="00:01:41.66" resultid="2584" heatid="4979" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="146" swimtime="00:00:47.35" resultid="2586" heatid="5130" lane="5" entrytime="00:00:54.26" entrycourse="SCM" />
                <RESULT eventid="4421" points="147" swimtime="00:00:41.16" resultid="5472" heatid="4761" lane="4" />
                <RESULT eventid="4445" points="143" swimtime="00:00:47.64" resultid="10316" heatid="6034" lane="6" />
                <RESULT eventid="10329" points="167" swimtime="00:00:36.59" resultid="10432" heatid="10345" lane="8" entrytime="00:00:36.86" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco" lastname="Crescente Rastelli" birthdate="2015-01-21" gender="M" nation="BRA" license="416673" swrid="5756904" athleteid="3059" externalid="416673" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" status="DNS" swimtime="00:00:00.00" resultid="3060" heatid="4751" lane="2" />
                <RESULT eventid="1102" status="DNS" swimtime="00:00:00.00" resultid="3061" heatid="4811" lane="2" />
                <RESULT eventid="1213" status="DNS" swimtime="00:00:00.00" resultid="3062" heatid="4951" lane="1" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="3063" heatid="4999" lane="1" />
                <RESULT eventid="1326" status="DNS" swimtime="00:00:00.00" resultid="3065" heatid="5126" lane="1" />
                <RESULT eventid="10329" status="DNS" swimtime="00:00:00.00" resultid="10466" heatid="10340" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="Pellanda" birthdate="2010-11-12" gender="M" nation="BRA" license="356352" swrid="5600233" athleteid="2183" externalid="356352" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="384" swimtime="00:00:29.90" resultid="2184" heatid="4773" lane="2" />
                <RESULT eventid="1105" points="331" swimtime="00:00:31.95" resultid="2185" heatid="4823" lane="5" />
                <RESULT eventid="1227" points="566" swimtime="00:02:00.08" resultid="2186" heatid="4965" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.00" />
                    <SPLIT distance="100" swimtime="00:00:58.17" />
                    <SPLIT distance="150" swimtime="00:01:28.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="484" swimtime="00:00:57.11" resultid="2187" heatid="5010" lane="4" entrytime="00:00:58.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="346" swimtime="00:00:35.51" resultid="2189" heatid="5140" lane="6" />
                <RESULT eventid="4423" points="384" swimtime="00:00:29.91" resultid="5540" heatid="4798" lane="3" />
                <RESULT eventid="4425" points="322" swimtime="00:00:31.70" resultid="5546" heatid="4807" lane="3" />
                <RESULT eventid="4429" points="324" swimtime="00:00:32.16" resultid="5577" heatid="4858" lane="2" />
                <RESULT eventid="4431" points="261" swimtime="00:00:34.59" resultid="5583" heatid="4867" lane="2" />
                <RESULT eventid="5807" points="380" swimtime="00:00:34.44" resultid="10287" heatid="6042" lane="3" />
                <RESULT eventid="10332" points="405" swimtime="00:00:27.24" resultid="10400" heatid="10357" lane="3" entrytime="00:00:28.13" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcelo" lastname="Luparia Vanhazebrock" birthdate="2010-01-31" gender="M" nation="BRA" athleteid="10339" externalid="339043" level="CLBO">
              <RESULTS>
                <RESULT eventid="10332" points="395" swimtime="00:00:27.46" resultid="10543" heatid="10346" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martina" lastname="Tallao Benke" birthdate="2012-01-02" gender="F" nation="BRA" license="376984" swrid="5588931" athleteid="2510" externalid="376984" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="527" swimtime="00:00:30.17" resultid="2511" heatid="4658" lane="6" />
                <RESULT eventid="1077" points="488" swimtime="00:00:32.05" resultid="2512" heatid="4722" lane="2" entrytime="00:00:34.22" entrycourse="SCM" />
                <RESULT eventid="1119" points="473" swimtime="00:02:32.63" resultid="2513" heatid="4876" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.78" />
                    <SPLIT distance="100" swimtime="00:01:13.71" />
                    <SPLIT distance="150" swimtime="00:01:54.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="456" swimtime="00:01:10.21" resultid="2514" heatid="4901" lane="4" entrytime="00:01:10.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="513" swimtime="00:00:28.63" resultid="2515" heatid="5097" lane="2" entrytime="00:00:28.55" entrycourse="SCM" />
                <RESULT eventid="1301" points="329" swimtime="00:00:41.09" resultid="2516" heatid="5034" lane="6" />
                <RESULT eventid="4411" points="498" swimtime="00:00:30.75" resultid="5387" heatid="4680" lane="1" />
                <RESULT eventid="4413" points="470" swimtime="00:00:31.35" resultid="5393" heatid="4691" lane="1" />
                <RESULT eventid="4417" points="466" swimtime="00:00:32.56" resultid="5417" heatid="4731" lane="1" />
                <RESULT eventid="4419" points="432" swimtime="00:00:33.39" resultid="5423" heatid="4742" lane="1" />
                <RESULT eventid="5801" points="342" swimtime="00:00:40.56" resultid="10102" heatid="6068" lane="6" />
                <RESULT eventid="5804" points="531" swimtime="00:00:28.31" resultid="10194" heatid="6054" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olivia" lastname="Mayer Paludetto" birthdate="2016-04-01" gender="F" nation="BRA" license="412014" swrid="5740014" athleteid="3025" externalid="412014" level="CLBO">
              <RESULTS>
                <RESULT eventid="1117" points="81" swimtime="00:00:58.14" resultid="3026" heatid="4872" lane="4" />
                <RESULT eventid="1141" points="104" swimtime="00:01:00.25" resultid="3027" heatid="4891" lane="4" />
                <RESULT eventid="1177" points="98" swimtime="00:00:49.70" resultid="3028" heatid="4918" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Fernandes Tramujas" birthdate="2015-01-15" gender="F" nation="BRA" license="406750" swrid="5717263" athleteid="2935" externalid="406750" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" status="DNS" swimtime="00:00:00.00" resultid="2936" heatid="4647" lane="5" entrytime="00:01:18.61" entrycourse="SCM" />
                <RESULT eventid="1074" status="DNS" swimtime="00:00:00.00" resultid="2937" heatid="4697" lane="3" entrytime="00:01:03.83" entrycourse="SCM" />
                <RESULT eventid="1129" status="DNS" swimtime="00:00:00.00" resultid="2938" heatid="4882" lane="1" />
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="2939" heatid="4909" lane="5" />
                <RESULT eventid="1298" status="DNS" swimtime="00:00:00.00" resultid="2940" heatid="5021" lane="6" entrytime="00:01:13.59" entrycourse="SCM" />
                <RESULT eventid="1311" status="DNS" swimtime="00:00:00.00" resultid="2941" heatid="5071" lane="5" entrytime="00:00:52.58" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Karam Barbosa Lima" birthdate="2012-12-11" gender="F" nation="BRA" license="376956" swrid="5588758" athleteid="2454" externalid="376956" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="276" swimtime="00:00:37.42" resultid="2455" heatid="4660" lane="5" />
                <RESULT eventid="1077" points="277" swimtime="00:00:38.70" resultid="2456" heatid="4720" lane="4" entrytime="00:00:37.51" entrycourse="SCM" />
                <RESULT eventid="1119" points="312" swimtime="00:02:55.26" resultid="2457" heatid="4875" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                    <SPLIT distance="100" swimtime="00:01:26.54" />
                    <SPLIT distance="150" swimtime="00:02:12.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="300" swimtime="00:01:21.91" resultid="2458" heatid="4913" lane="4" entrytime="00:01:22.38" entrycourse="SCM" />
                <RESULT eventid="1314" points="323" swimtime="00:00:33.41" resultid="2459" heatid="5093" lane="6" entrytime="00:00:32.38" entrycourse="SCM" />
                <RESULT eventid="1301" points="228" swimtime="00:00:46.38" resultid="2460" heatid="5037" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giuliana" lastname="Sovierzoski Ferreira" birthdate="2015-01-20" gender="F" nation="BRA" license="397168" swrid="5641776" athleteid="2809" externalid="397168" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" status="DNS" swimtime="00:00:00.00" resultid="2810" heatid="4647" lane="1" entrytime="00:01:19.82" entrycourse="SCM" />
                <RESULT eventid="1074" status="DNS" swimtime="00:00:00.00" resultid="2811" heatid="4698" lane="3" entrytime="00:00:56.97" entrycourse="SCM" />
                <RESULT eventid="1129" points="162" swimtime="00:01:54.16" resultid="2812" heatid="4883" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="91" swimtime="00:02:01.94" resultid="2813" heatid="4905" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="152" swimtime="00:00:53.15" resultid="2814" heatid="5025" lane="7" entrytime="00:00:53.07" entrycourse="SCM" />
                <RESULT eventid="1311" points="127" swimtime="00:00:45.54" resultid="2815" heatid="5072" lane="1" entrytime="00:00:50.08" entrycourse="SCM" />
                <RESULT eventid="4433" points="159" swimtime="00:00:52.33" resultid="10083" heatid="5029" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Della Villa Yang" birthdate="2015-02-27" gender="F" nation="BRA" license="393283" swrid="5616442" athleteid="2788" externalid="393283" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="176" swimtime="00:00:43.46" resultid="2789" heatid="4651" lane="6" entrytime="00:00:46.47" entrycourse="SCM" />
                <RESULT eventid="1074" points="158" swimtime="00:00:46.69" resultid="2790" heatid="4701" lane="6" entrytime="00:00:49.19" entrycourse="SCM" />
                <RESULT eventid="1129" points="170" swimtime="00:01:52.48" resultid="2791" heatid="4880" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="115" swimtime="00:01:51.08" resultid="2792" heatid="4898" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="165" swimtime="00:00:51.64" resultid="2793" heatid="5023" lane="7" entrytime="00:01:02.88" entrycourse="SCM" />
                <RESULT eventid="1311" points="206" swimtime="00:00:38.78" resultid="2794" heatid="5075" lane="4" entrytime="00:00:40.03" entrycourse="SCM" />
                <RESULT eventid="4409" points="157" swimtime="00:00:45.10" resultid="5363" heatid="4655" lane="1" />
                <RESULT eventid="4415" points="148" swimtime="00:00:47.66" resultid="5400" heatid="4706" lane="5" />
                <RESULT eventid="4433" points="163" swimtime="00:00:51.88" resultid="10082" heatid="5029" lane="4" />
                <RESULT eventid="4439" points="201" swimtime="00:00:39.08" resultid="10175" heatid="6048" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="De Lima Cavalcanti" birthdate="2014-10-07" gender="M" nation="BRA" license="385884" swrid="5684550" athleteid="2879" externalid="385884" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="122" swimtime="00:00:43.82" resultid="2880" heatid="4755" lane="3" entrytime="00:00:43.98" entrycourse="SCM" />
                <RESULT eventid="1102" points="159" swimtime="00:00:40.75" resultid="2881" heatid="4817" lane="4" entrytime="00:00:40.24" entrycourse="SCM" />
                <RESULT eventid="1249" points="171" swimtime="00:01:27.07" resultid="2882" heatid="4983" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1237" points="101" swimtime="00:01:42.48" resultid="2883" heatid="4969" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="113" swimtime="00:00:51.49" resultid="2885" heatid="5124" lane="5" />
                <RESULT eventid="4427" points="169" swimtime="00:00:39.99" resultid="5507" heatid="4822" lane="3" />
                <RESULT eventid="10329" points="180" swimtime="00:00:35.66" resultid="10450" heatid="10344" lane="5" entrytime="00:00:37.61" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Albuquerque" birthdate="2012-08-17" gender="F" nation="BRA" license="369275" swrid="5602507" athleteid="2370" externalid="369275" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="288" swimtime="00:00:36.89" resultid="2371" heatid="4670" lane="2" entrytime="00:00:36.53" entrycourse="SCM" />
                <RESULT eventid="1077" points="216" swimtime="00:00:42.02" resultid="2372" heatid="4709" lane="2" />
                <RESULT eventid="1129" points="439" swimtime="00:01:22.02" resultid="2373" heatid="4887" lane="5" entrytime="00:01:22.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="407" swimtime="00:03:01.58" resultid="2374" heatid="4921" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.28" />
                    <SPLIT distance="100" swimtime="00:01:26.75" />
                    <SPLIT distance="150" swimtime="00:02:15.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="303" swimtime="00:00:34.12" resultid="2375" heatid="5092" lane="1" entrytime="00:00:33.16" entrycourse="SCM" />
                <RESULT eventid="1301" points="393" swimtime="00:00:38.73" resultid="2376" heatid="5045" lane="5" entrytime="00:00:37.52" entrycourse="SCM" />
                <RESULT eventid="5801" points="401" swimtime="00:00:38.46" resultid="10097" heatid="6068" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Saber" birthdate="2014-06-04" gender="F" nation="BRA" license="392141" swrid="5602554" athleteid="2732" externalid="392141" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="88" swimtime="00:00:54.64" resultid="2733" heatid="4649" lane="6" entrytime="00:00:56.24" entrycourse="SCM" />
                <RESULT eventid="1074" points="135" swimtime="00:00:49.20" resultid="2734" heatid="4701" lane="2" entrytime="00:00:48.59" entrycourse="SCM" />
                <RESULT eventid="1129" points="215" swimtime="00:01:44.09" resultid="2735" heatid="4881" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:44.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="131" swimtime="00:01:48.05" resultid="2736" heatid="4906" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="196" swimtime="00:00:48.82" resultid="2737" heatid="5025" lane="5" entrytime="00:00:50.06" entrycourse="SCM" />
                <RESULT eventid="1311" points="187" swimtime="00:00:40.07" resultid="2738" heatid="5075" lane="8" entrytime="00:00:42.37" entrycourse="SCM" />
                <RESULT eventid="4433" points="190" swimtime="00:00:49.27" resultid="10089" heatid="6064" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Ribas Luz" birthdate="2015-02-05" gender="F" nation="BRA" license="406743" swrid="5717291" athleteid="2900" externalid="406743" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="52" swimtime="00:01:05.22" resultid="2901" heatid="4646" lane="3" entrytime="00:01:37.59" entrycourse="SCM" />
                <RESULT eventid="1074" points="93" swimtime="00:00:55.63" resultid="2902" heatid="4699" lane="2" entrytime="00:00:54.00" entrycourse="SCM" />
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="2903" heatid="4909" lane="4" />
                <RESULT eventid="1189" status="DNS" swimtime="00:00:00.00" resultid="2904" heatid="4926" lane="4" entrytime="00:02:03.43" entrycourse="SCM" />
                <RESULT eventid="1298" status="DNS" swimtime="00:00:00.00" resultid="2905" heatid="5021" lane="2" entrytime="00:01:08.95" entrycourse="SCM" />
                <RESULT eventid="1311" status="DNS" swimtime="00:00:00.00" resultid="2906" heatid="5071" lane="1" entrytime="00:00:55.24" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Pisani Ferreira" birthdate="2014-01-26" gender="M" nation="BRA" license="391017" swrid="5602570" athleteid="2648" externalid="391017" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" status="DNS" swimtime="00:00:00.00" resultid="2649" heatid="4754" lane="1" entrytime="00:00:54.17" entrycourse="SCM" />
                <RESULT eventid="1102" status="DNS" swimtime="00:00:00.00" resultid="2650" heatid="4811" lane="1" />
                <RESULT eventid="1213" status="DNS" swimtime="00:00:00.00" resultid="2651" heatid="4948" lane="3" />
                <RESULT eventid="1249" status="DNS" swimtime="00:00:00.00" resultid="2652" heatid="4978" lane="4" />
                <RESULT eventid="1326" status="DNS" swimtime="00:00:00.00" resultid="2654" heatid="5131" lane="1" entrytime="00:00:50.93" entrycourse="SCM" />
                <RESULT eventid="10329" status="DNS" swimtime="00:00:00.00" resultid="10438" heatid="10343" lane="6" entrytime="00:00:41.70" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Da Cunha Souza" birthdate="2015-05-30" gender="F" nation="BRA" license="400016" swrid="5652883" athleteid="2844" externalid="400016" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="132" swimtime="00:00:47.77" resultid="2845" heatid="4649" lane="5" entrytime="00:00:54.69" entrycourse="SCM" />
                <RESULT eventid="1074" points="170" swimtime="00:00:45.53" resultid="2846" heatid="4701" lane="4" entrytime="00:00:48.55" entrycourse="SCM" />
                <RESULT eventid="1165" points="161" swimtime="00:01:40.74" resultid="2847" heatid="4905" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="174" swimtime="00:01:29.96" resultid="2848" heatid="4927" lane="5" entrytime="00:01:37.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="115" swimtime="00:00:58.24" resultid="2849" heatid="5023" lane="6" entrytime="00:01:02.80" entrycourse="SCM" />
                <RESULT eventid="1311" points="238" swimtime="00:00:36.96" resultid="2850" heatid="5075" lane="2" entrytime="00:00:40.69" entrycourse="SCM" />
                <RESULT eventid="4409" points="134" swimtime="00:00:47.62" resultid="5366" heatid="4655" lane="4" />
                <RESULT eventid="4415" points="171" swimtime="00:00:45.46" resultid="5397" heatid="4706" lane="2" />
                <RESULT eventid="4433" points="132" swimtime="00:00:55.66" resultid="10078" heatid="5029" lane="1" />
                <RESULT eventid="4439" points="250" swimtime="00:00:36.37" resultid="10174" heatid="6048" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Menezes" birthdate="2015-07-28" gender="F" nation="BRA" license="412898" swrid="5755339" athleteid="3040" externalid="412898" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="40" swimtime="00:01:11.07" resultid="3041" heatid="4646" lane="2" />
                <RESULT eventid="1074" points="110" swimtime="00:00:52.64" resultid="3042" heatid="4696" lane="1" />
                <RESULT eventid="1165" points="106" swimtime="00:01:55.65" resultid="3043" heatid="4906" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="103" swimtime="00:01:47.07" resultid="3044" heatid="4925" lane="4" />
                <RESULT eventid="1298" status="DNS" swimtime="00:00:00.00" resultid="3045" heatid="5020" lane="2" />
                <RESULT eventid="1311" points="133" swimtime="00:00:44.85" resultid="3046" heatid="5071" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Rocha" birthdate="2011-08-25" gender="F" nation="BRA" license="366904" swrid="5602578" athleteid="2281" externalid="366904" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="395" swimtime="00:00:33.21" resultid="2282" heatid="4664" lane="6" />
                <RESULT eventid="1077" points="320" swimtime="00:00:36.89" resultid="2283" heatid="4710" lane="2" />
                <RESULT eventid="1119" points="380" swimtime="00:02:44.16" resultid="2284" heatid="4875" lane="6" />
                <RESULT eventid="1153" points="291" swimtime="00:01:21.56" resultid="2285" heatid="4899" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="417" swimtime="00:00:30.68" resultid="2286" heatid="5084" lane="2" />
                <RESULT eventid="1301" points="264" swimtime="00:00:44.19" resultid="2287" heatid="5036" lane="3" />
                <RESULT eventid="4411" points="398" swimtime="00:00:33.13" resultid="5353" heatid="4682" lane="1" />
                <RESULT eventid="4413" points="403" swimtime="00:00:32.98" resultid="5359" heatid="4692" lane="1" />
                <RESULT eventid="4417" points="331" swimtime="00:00:36.47" resultid="5430" heatid="4733" lane="5" />
                <RESULT eventid="5804" points="432" swimtime="00:00:30.33" resultid="10201" heatid="6056" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Poletto Abrahao" birthdate="2014-10-20" gender="M" nation="BRA" license="382128" swrid="5602571" athleteid="2594" externalid="382128" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="181" swimtime="00:00:38.40" resultid="2595" heatid="4756" lane="4" entrytime="00:00:39.22" entrycourse="SCM" />
                <RESULT eventid="1102" points="125" swimtime="00:00:44.14" resultid="2596" heatid="4812" lane="6" />
                <RESULT eventid="1213" points="188" swimtime="00:01:36.44" resultid="2597" heatid="4951" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="136" swimtime="00:01:33.88" resultid="2598" heatid="4980" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="196" swimtime="00:00:42.92" resultid="2600" heatid="5131" lane="3" entrytime="00:00:42.87" entrycourse="SCM" />
                <RESULT eventid="4421" points="164" swimtime="00:00:39.70" resultid="5470" heatid="4761" lane="2" />
                <RESULT eventid="4427" points="136" swimtime="00:00:42.92" resultid="5509" heatid="4822" lane="5" />
                <RESULT eventid="4445" points="204" swimtime="00:00:42.33" resultid="10314" heatid="6034" lane="4" />
                <RESULT eventid="10329" points="203" swimtime="00:00:34.29" resultid="10434" heatid="10345" lane="5" entrytime="00:00:35.36" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Alice Palhano" birthdate="2016-04-06" gender="F" nation="BRA" license="412015" swrid="5740004" athleteid="3029" externalid="412015" level="CLBO">
              <RESULTS>
                <RESULT eventid="1117" points="46" swimtime="00:01:10.07" resultid="3030" heatid="4872" lane="2" />
                <RESULT eventid="1141" points="54" swimtime="00:01:14.70" resultid="3031" heatid="4891" lane="2" />
                <RESULT eventid="1177" points="39" swimtime="00:01:07.29" resultid="3032" heatid="4918" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Antunes Saboia" birthdate="2012-06-28" gender="M" nation="BRA" license="369278" swrid="5602511" athleteid="2391" externalid="369278" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="185" swimtime="00:00:38.14" resultid="2392" heatid="4767" lane="1" />
                <RESULT eventid="1105" points="189" swimtime="00:00:38.48" resultid="2393" heatid="4836" lane="1" entrytime="00:00:41.34" entrycourse="SCM" />
                <RESULT eventid="1213" points="271" swimtime="00:01:25.38" resultid="2394" heatid="4953" lane="1" entrytime="00:01:27.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="282" swimtime="00:03:03.23" resultid="2395" heatid="4992" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.08" />
                    <SPLIT distance="100" swimtime="00:01:30.45" />
                    <SPLIT distance="150" swimtime="00:02:17.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="270" swimtime="00:00:38.56" resultid="2397" heatid="5152" lane="8" entrytime="00:00:39.02" entrycourse="SCM" />
                <RESULT eventid="5807" points="267" swimtime="00:00:38.74" resultid="10277" heatid="6038" lane="6" />
                <RESULT eventid="10332" points="269" swimtime="00:00:31.23" resultid="10418" heatid="10353" lane="1" entrytime="00:00:32.56" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Magalhaes Dos Reis" birthdate="2010-05-05" gender="M" nation="BRA" license="356361" swrid="5600207" athleteid="2225" externalid="356361" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="387" swimtime="00:00:29.83" resultid="2226" heatid="4768" lane="4" />
                <RESULT eventid="1105" points="205" swimtime="00:00:37.44" resultid="2227" heatid="5253" lane="2" />
                <RESULT eventid="1237" points="299" swimtime="00:01:11.40" resultid="2228" heatid="4973" lane="5" entrytime="00:01:15.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="378" swimtime="00:01:01.98" resultid="2229" heatid="5010" lane="6" entrytime="00:01:00.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="286" swimtime="00:00:37.84" resultid="2231" heatid="5139" lane="6" />
                <RESULT eventid="4423" points="369" swimtime="00:00:30.31" resultid="5539" heatid="4798" lane="2" />
                <RESULT eventid="10332" points="399" swimtime="00:00:27.38" resultid="10404" heatid="10358" lane="2" entrytime="00:00:27.78" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Liam" lastname="Batista Grise" birthdate="2014-03-27" gender="M" nation="BRA" license="391008" swrid="5602514" athleteid="2629" externalid="391008" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" status="DNS" swimtime="00:00:00.00" resultid="2630" heatid="4752" lane="5" />
                <RESULT eventid="1102" status="DNS" swimtime="00:00:00.00" resultid="2631" heatid="4815" lane="6" entrytime="00:00:52.62" entrycourse="SCM" />
                <RESULT eventid="1213" status="DNS" swimtime="00:00:00.00" resultid="2632" heatid="4949" lane="3" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="2633" heatid="5002" lane="6" entrytime="00:01:43.32" entrycourse="SCM" />
                <RESULT eventid="1326" status="DNS" swimtime="00:00:00.00" resultid="2635" heatid="5130" lane="4" entrytime="00:00:53.14" entrycourse="SCM" />
                <RESULT eventid="10329" status="DNS" swimtime="00:00:00.00" resultid="10437" heatid="10343" lane="5" entrytime="00:00:40.55" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Coelho Ghignone" birthdate="2015-01-05" gender="M" nation="BRA" license="410201" swrid="5740006" athleteid="3011" externalid="410201" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="128" swimtime="00:00:43.12" resultid="3012" heatid="4749" lane="2" />
                <RESULT eventid="1102" points="128" swimtime="00:00:43.81" resultid="3013" heatid="4815" lane="4" entrytime="00:00:50.09" entrycourse="SCM" />
                <RESULT eventid="1249" status="DNS" swimtime="00:00:00.00" resultid="3014" heatid="4979" lane="5" />
                <RESULT eventid="1273" points="159" swimtime="00:01:22.73" resultid="3015" heatid="5002" lane="2" entrytime="00:01:37.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="101" swimtime="00:00:53.53" resultid="3017" heatid="5128" lane="6" entrytime="00:01:05.25" entrycourse="SCM" />
                <RESULT eventid="4421" points="129" swimtime="00:00:43.02" resultid="5465" heatid="4760" lane="3" />
                <RESULT eventid="4427" points="132" swimtime="00:00:43.32" resultid="5500" heatid="4821" lane="2" />
                <RESULT eventid="4445" points="100" swimtime="00:00:53.61" resultid="10306" heatid="6032" lane="2" />
                <RESULT eventid="10329" points="166" swimtime="00:00:36.66" resultid="10461" heatid="10343" lane="1" entrytime="00:00:40.89" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Barbara" lastname="Bittencourt Ribas" birthdate="2013-02-01" gender="F" nation="BRA" license="372682" swrid="5588555" athleteid="2433" externalid="372682" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="269" swimtime="00:00:37.76" resultid="2434" heatid="4668" lane="2" entrytime="00:00:39.28" entrycourse="SCM" />
                <RESULT eventid="1077" points="269" swimtime="00:00:39.11" resultid="2435" heatid="4717" lane="4" entrytime="00:00:41.60" entrycourse="SCM" />
                <RESULT eventid="1119" points="321" swimtime="00:02:53.57" resultid="2436" heatid="4875" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                    <SPLIT distance="100" swimtime="00:01:27.03" />
                    <SPLIT distance="150" swimtime="00:02:12.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="310" swimtime="00:01:21.10" resultid="2437" heatid="4913" lane="2" entrytime="00:01:23.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="348" swimtime="00:00:32.59" resultid="2438" heatid="5090" lane="7" entrytime="00:00:33.28" entrycourse="SCM" />
                <RESULT eventid="1301" status="DNS" swimtime="00:00:00.00" resultid="2439" heatid="5040" lane="2" entrytime="00:00:48.97" entrycourse="SCM" />
                <RESULT eventid="4417" points="283" swimtime="00:00:38.43" resultid="5410" heatid="4729" lane="3" />
                <RESULT eventid="4419" points="289" swimtime="00:00:38.17" resultid="5416" heatid="4741" lane="3" />
                <RESULT eventid="5804" points="324" swimtime="00:00:33.38" resultid="10191" heatid="6052" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Brandt Macedo" birthdate="2013-04-19" gender="M" nation="BRA" license="414421" swrid="5755329" athleteid="3054" externalid="414421" level="CLBO">
              <RESULTS>
                <RESULT comment="SW 8.3 - Movimento alternado das pernas ou pés., SW 8.3 - Movimento de pernada de peito." eventid="1092" status="DSQ" swimtime="00:01:12.38" resultid="3055" heatid="4770" lane="1" />
                <RESULT comment="SW 6.5 - Não terminou a prova enquanto estava de costas.&#10;&#10;&#10;&#10;&#10;&#10;&#10;" eventid="1105" status="DSQ" swimtime="00:01:06.83" resultid="3056" heatid="4828" lane="5" />
                <RESULT eventid="1329" points="88" swimtime="00:00:56.07" resultid="3058" heatid="5143" lane="4" />
                <RESULT eventid="10332" points="47" swimtime="00:00:55.79" resultid="10465" heatid="10347" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniela" lastname="Dolberth Alcantara" birthdate="2014-09-26" gender="F" nation="BRA" license="382124" swrid="5602532" athleteid="2573" externalid="382124" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="154" swimtime="00:00:45.44" resultid="2574" heatid="4650" lane="1" entrytime="00:00:51.49" entrycourse="SCM" />
                <RESULT eventid="1074" points="166" swimtime="00:00:45.91" resultid="2575" heatid="4700" lane="5" entrytime="00:00:51.72" entrycourse="SCM" />
                <RESULT eventid="1129" points="158" swimtime="00:01:55.25" resultid="2576" heatid="4882" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="162" swimtime="00:01:40.69" resultid="2577" heatid="4910" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="141" swimtime="00:00:54.44" resultid="2578" heatid="5024" lane="8" entrytime="00:00:57.72" entrycourse="SCM" />
                <RESULT eventid="1311" points="194" swimtime="00:00:39.57" resultid="2579" heatid="5073" lane="1" entrytime="00:00:44.38" entrycourse="SCM" />
                <RESULT eventid="4409" points="173" swimtime="00:00:43.70" resultid="5374" heatid="4656" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enrico" lastname="Hallage Bianchini" birthdate="2014-02-27" gender="M" nation="BRA" license="397164" swrid="5661348" athleteid="2802" externalid="397164" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" status="DNS" swimtime="00:00:00.00" resultid="2803" heatid="4756" lane="1" entrytime="00:00:43.35" entrycourse="SCM" />
                <RESULT eventid="1102" status="DNS" swimtime="00:00:00.00" resultid="2804" heatid="4816" lane="2" entrytime="00:00:44.70" entrycourse="SCM" />
                <RESULT eventid="1249" status="DNS" swimtime="00:00:00.00" resultid="2805" heatid="4978" lane="1" />
                <RESULT eventid="1237" status="DNS" swimtime="00:00:00.00" resultid="2806" heatid="4969" lane="2" />
                <RESULT eventid="1326" status="DNS" swimtime="00:00:00.00" resultid="2808" heatid="5124" lane="6" />
                <RESULT eventid="10329" status="DNS" swimtime="00:00:00.00" resultid="10447" heatid="10344" lane="8" entrytime="00:00:39.66" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Gois Nogueira" birthdate="2014-03-11" gender="F" nation="BRA" license="393258" swrid="5616443" athleteid="2739" externalid="393258" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="83" swimtime="00:00:55.87" resultid="2740" heatid="4650" lane="6" entrytime="00:00:52.11" entrycourse="SCM" />
                <RESULT eventid="1074" points="136" swimtime="00:00:49.02" resultid="2741" heatid="4700" lane="3" entrytime="00:00:49.71" entrycourse="SCM" />
                <RESULT eventid="1129" points="157" swimtime="00:01:55.43" resultid="2742" heatid="4883" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="125" swimtime="00:01:49.49" resultid="2743" heatid="4907" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="175" swimtime="00:00:50.66" resultid="2744" heatid="5024" lane="3" entrytime="00:00:53.12" entrycourse="SCM" />
                <RESULT eventid="1311" points="203" swimtime="00:00:38.96" resultid="2745" heatid="5075" lane="3" entrytime="00:00:39.64" entrycourse="SCM" />
                <RESULT eventid="4433" points="208" swimtime="00:00:47.85" resultid="10090" heatid="6064" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Leao" birthdate="2011-09-18" gender="M" nation="BRA" license="366880" swrid="5602553" athleteid="2232" externalid="366880" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="300" swimtime="00:00:32.49" resultid="2233" heatid="4762" lane="3" />
                <RESULT eventid="1105" points="250" swimtime="00:00:35.07" resultid="2234" heatid="4824" lane="4" />
                <RESULT eventid="1227" points="387" swimtime="00:02:16.26" resultid="2235" heatid="4965" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:06.98" />
                    <SPLIT distance="150" swimtime="00:01:42.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="363" swimtime="00:01:02.81" resultid="2236" heatid="4999" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="221" swimtime="00:00:41.23" resultid="2238" heatid="5140" lane="4" />
                <RESULT eventid="10332" points="351" swimtime="00:00:28.57" resultid="10405" heatid="10356" lane="3" entrytime="00:00:29.57" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="LIV" lastname="Carvalho" birthdate="2011-09-13" gender="F" nation="BRA" license="366899" swrid="5602524" athleteid="2267" externalid="366899" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="254" swimtime="00:00:38.48" resultid="2268" heatid="4661" lane="3" />
                <RESULT eventid="1077" points="175" swimtime="00:00:45.14" resultid="2269" heatid="4709" lane="5" />
                <RESULT eventid="1129" points="342" swimtime="00:01:29.12" resultid="2270" heatid="4885" lane="2" entrytime="00:01:36.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="311" swimtime="00:01:14.13" resultid="2271" heatid="4929" lane="3" entrytime="00:01:17.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="308" swimtime="00:00:33.95" resultid="2272" heatid="5083" lane="4" />
                <RESULT eventid="1301" points="338" swimtime="00:00:40.69" resultid="2273" heatid="5036" lane="6" />
                <RESULT eventid="5801" points="342" swimtime="00:00:40.55" resultid="10157" heatid="6070" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Szpak Zraik" birthdate="2015-04-10" gender="M" nation="BRA" license="393259" swrid="5616451" athleteid="2746" externalid="393259" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="109" swimtime="00:00:45.52" resultid="2747" heatid="4754" lane="3" entrytime="00:00:49.44" entrycourse="SCM" />
                <RESULT eventid="1102" points="94" swimtime="00:00:48.46" resultid="2748" heatid="4811" lane="3" />
                <RESULT eventid="1213" points="163" swimtime="00:01:41.08" resultid="2749" heatid="4950" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="82" swimtime="00:01:51.04" resultid="2750" heatid="4982" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="158" swimtime="00:00:46.13" resultid="2752" heatid="5131" lane="4" entrytime="00:00:48.08" entrycourse="SCM" />
                <RESULT eventid="4421" points="116" swimtime="00:00:44.53" resultid="5466" heatid="4760" lane="4" />
                <RESULT eventid="4445" points="164" swimtime="00:00:45.49" resultid="10308" heatid="6032" lane="4" />
                <RESULT eventid="4427" points="93" swimtime="00:00:48.79" resultid="10326" heatid="4821" lane="6" />
                <RESULT eventid="10329" points="126" swimtime="00:00:40.20" resultid="10444" heatid="10344" lane="7" entrytime="00:00:39.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Magalhaes Dabul" birthdate="2014-01-05" gender="M" nation="BRA" license="391023" swrid="5602555" athleteid="2683" externalid="391023" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="135" swimtime="00:00:42.38" resultid="2684" heatid="4755" lane="4" entrytime="00:00:44.09" entrycourse="SCM" />
                <RESULT eventid="1102" points="99" swimtime="00:00:47.70" resultid="2685" heatid="4814" lane="5" entrytime="00:00:55.28" entrycourse="SCM" />
                <RESULT eventid="1213" points="145" swimtime="00:01:45.00" resultid="2686" heatid="4949" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1237" points="103" swimtime="00:01:41.90" resultid="2687" heatid="4971" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="141" swimtime="00:00:47.85" resultid="2689" heatid="5124" lane="2" />
                <RESULT eventid="4421" points="139" swimtime="00:00:41.91" resultid="5473" heatid="4761" lane="5" />
                <RESULT eventid="4445" points="150" swimtime="00:00:46.92" resultid="10312" heatid="6034" lane="2" />
                <RESULT eventid="10329" points="157" swimtime="00:00:37.30" resultid="10441" heatid="10345" lane="7" entrytime="00:00:37.78" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Bernardi Pedrosa" birthdate="2013-03-09" gender="F" nation="BRA" license="376977" swrid="5588551" athleteid="2496" externalid="376977" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="177" swimtime="00:00:43.36" resultid="2497" heatid="4660" lane="6" />
                <RESULT eventid="1077" points="264" swimtime="00:00:39.36" resultid="2498" heatid="4719" lane="5" entrytime="00:00:39.52" entrycourse="SCM" />
                <RESULT eventid="1119" points="271" swimtime="00:03:03.66" resultid="2499" heatid="4875" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.22" />
                    <SPLIT distance="100" swimtime="00:01:31.50" />
                    <SPLIT distance="150" swimtime="00:02:19.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="250" swimtime="00:01:27.13" resultid="2500" heatid="4913" lane="6" entrytime="00:01:28.68" entrycourse="SCM" />
                <RESULT eventid="1314" points="288" swimtime="00:00:34.71" resultid="2501" heatid="5089" lane="2" entrytime="00:00:35.23" entrycourse="SCM" />
                <RESULT eventid="1301" points="178" swimtime="00:00:50.42" resultid="2502" heatid="5037" lane="4" />
                <RESULT eventid="4417" points="252" swimtime="00:00:39.97" resultid="5411" heatid="4729" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elisa" lastname="Osternack Almeida" birthdate="2015-04-14" gender="F" nation="BRA" license="406747" swrid="5717286" athleteid="2914" externalid="406747" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" status="DNS" swimtime="00:00:00.00" resultid="2915" heatid="4648" lane="2" entrytime="00:00:59.52" entrycourse="SCM" />
                <RESULT eventid="1074" status="DNS" swimtime="00:00:00.00" resultid="2916" heatid="4699" lane="3" entrytime="00:00:53.12" entrycourse="SCM" />
                <RESULT eventid="1129" status="DNS" swimtime="00:00:00.00" resultid="2917" heatid="4880" lane="4" />
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="2918" heatid="4909" lane="6" />
                <RESULT eventid="1298" status="DNS" swimtime="00:00:00.00" resultid="2919" heatid="5020" lane="4" />
                <RESULT eventid="1311" status="DNS" swimtime="00:00:00.00" resultid="2920" heatid="5072" lane="2" entrytime="00:00:47.03" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Pens Correa" birthdate="2015-11-27" gender="M" nation="BRA" license="393262" swrid="5616449" athleteid="2767" externalid="393262" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="178" swimtime="00:00:38.63" resultid="2768" heatid="4756" lane="3" entrytime="00:00:38.61" entrycourse="SCM" />
                <RESULT eventid="1102" points="160" swimtime="00:00:40.67" resultid="2769" heatid="4817" lane="3" entrytime="00:00:39.23" entrycourse="SCM" />
                <RESULT eventid="1249" points="142" swimtime="00:01:32.56" resultid="2770" heatid="4983" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1237" points="127" swimtime="00:01:35.04" resultid="2771" heatid="4970" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="138" swimtime="00:00:48.18" resultid="2773" heatid="5124" lane="4" />
                <RESULT eventid="4421" points="182" swimtime="00:00:38.34" resultid="5463" heatid="4760" lane="1" />
                <RESULT eventid="4427" points="180" swimtime="00:00:39.15" resultid="5499" heatid="4821" lane="1" />
                <RESULT eventid="4445" points="142" swimtime="00:00:47.75" resultid="10307" heatid="6032" lane="3" />
                <RESULT eventid="10329" points="212" swimtime="00:00:33.80" resultid="10445" heatid="10345" lane="2" entrytime="00:00:34.98" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Guilherme Garcia" birthdate="2015-10-26" gender="M" nation="BRA" license="406967" swrid="5717271" athleteid="2990" externalid="406967" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" status="DNS" swimtime="00:00:00.00" resultid="2991" heatid="4753" lane="1" entrytime="00:01:29.25" entrycourse="SCM" />
                <RESULT eventid="1102" status="DNS" swimtime="00:00:00.00" resultid="2992" heatid="4812" lane="4" entrytime="00:01:04.75" entrycourse="SCM" />
                <RESULT eventid="1249" status="DNS" swimtime="00:00:00.00" resultid="2993" heatid="4978" lane="3" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="2994" heatid="5001" lane="1" entrytime="00:02:14.17" entrycourse="SCM" />
                <RESULT eventid="1326" status="DNS" swimtime="00:00:00.00" resultid="2996" heatid="5127" lane="6" entrytime="00:01:30.86" entrycourse="SCM" />
                <RESULT eventid="10329" status="DNS" swimtime="00:00:00.00" resultid="10460" heatid="10340" lane="3" entrytime="00:00:57.09" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Viera Correa" birthdate="2012-03-07" gender="M" nation="BRA" license="369269" swrid="5602590" athleteid="2344" externalid="369269" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="262" swimtime="00:00:33.98" resultid="2345" heatid="4777" lane="5" entrytime="00:00:37.05" entrycourse="SCM" />
                <RESULT eventid="1105" points="226" swimtime="00:00:36.29" resultid="2346" heatid="4837" lane="4" entrytime="00:00:38.50" entrycourse="SCM" />
                <RESULT eventid="1227" points="314" swimtime="00:02:26.09" resultid="2347" heatid="4966" lane="3" entrytime="00:02:38.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                    <SPLIT distance="100" swimtime="00:01:11.23" />
                    <SPLIT distance="150" swimtime="00:01:50.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="303" swimtime="00:01:06.70" resultid="2348" heatid="5007" lane="4" entrytime="00:01:06.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="200" swimtime="00:00:42.66" resultid="2350" heatid="5147" lane="6" />
                <RESULT eventid="4423" points="264" swimtime="00:00:33.90" resultid="5494" heatid="4794" lane="2" />
                <RESULT eventid="4429" points="230" swimtime="00:00:36.05" resultid="5523" heatid="4854" lane="4" />
                <RESULT eventid="4431" points="208" swimtime="00:00:37.29" resultid="5527" heatid="4865" lane="2" />
                <RESULT eventid="4425" points="209" swimtime="00:00:36.65" resultid="5604" heatid="4805" lane="2" />
                <RESULT eventid="10332" points="314" swimtime="00:00:29.64" resultid="10414" heatid="10355" lane="8" entrytime="00:00:30.32" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Simioni Albuquerque" birthdate="2014-12-23" gender="F" nation="BRA" license="401980" swrid="5661355" athleteid="2858" externalid="401980" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="240" swimtime="00:00:39.23" resultid="2859" heatid="4651" lane="4" entrytime="00:00:40.27" entrycourse="SCM" />
                <RESULT eventid="1074" points="185" swimtime="00:00:44.28" resultid="2860" heatid="4701" lane="5" entrytime="00:00:48.84" entrycourse="SCM" />
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente., Na chegada." eventid="1153" status="DSQ" swimtime="00:01:43.18" resultid="2861" heatid="4899" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="226" swimtime="00:01:22.45" resultid="2862" heatid="4927" lane="3" entrytime="00:01:33.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="204" swimtime="00:00:48.15" resultid="2863" heatid="5020" lane="6" />
                <RESULT eventid="1311" points="290" swimtime="00:00:34.62" resultid="2864" heatid="5076" lane="5" entrytime="00:00:37.22" entrycourse="SCM" />
                <RESULT eventid="4415" points="191" swimtime="00:00:43.81" resultid="5407" heatid="4707" lane="6" />
                <RESULT eventid="4433" points="197" swimtime="00:00:48.75" resultid="10088" heatid="6064" lane="4" />
                <RESULT eventid="4439" points="272" swimtime="00:00:35.39" resultid="10183" heatid="6050" lane="4" />
                <RESULT eventid="4409" points="206" swimtime="00:00:41.24" resultid="10323" heatid="4656" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Schiavo Vianna" birthdate="2013-04-27" gender="F" nation="BRA" license="391005" swrid="5602582" athleteid="2615" externalid="391005" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="93" swimtime="00:00:53.80" resultid="2616" heatid="4666" lane="5" entrytime="00:00:55.93" entrycourse="SCM" />
                <RESULT eventid="1077" points="154" swimtime="00:00:47.04" resultid="2617" heatid="4711" lane="1" />
                <RESULT eventid="1143" points="227" swimtime="00:03:00.59" resultid="2618" heatid="4894" lane="5" entrytime="00:03:33.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.41" />
                    <SPLIT distance="100" swimtime="00:01:25.22" />
                    <SPLIT distance="150" swimtime="00:02:12.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="228" swimtime="00:01:22.17" resultid="2619" heatid="4928" lane="2" entrytime="00:01:25.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="285" swimtime="00:00:34.84" resultid="2620" heatid="5086" lane="8" entrytime="00:00:36.82" entrycourse="SCM" />
                <RESULT eventid="1301" points="255" swimtime="00:00:44.72" resultid="2621" heatid="5040" lane="3" entrytime="00:00:48.50" entrycourse="SCM" />
                <RESULT eventid="5801" points="254" swimtime="00:00:44.76" resultid="10096" heatid="6066" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Afonso Fowler" birthdate="2014-01-22" gender="M" nation="BRA" license="393264" swrid="5661338" athleteid="2781" externalid="393264" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" status="DNS" swimtime="00:00:00.00" resultid="2782" heatid="4754" lane="6" entrytime="00:00:58.54" entrycourse="SCM" />
                <RESULT eventid="1102" status="DNS" swimtime="00:00:00.00" resultid="2783" heatid="4814" lane="4" entrytime="00:00:53.27" entrycourse="SCM" />
                <RESULT eventid="1249" status="DNS" swimtime="00:00:00.00" resultid="2784" heatid="4978" lane="6" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="2785" heatid="5003" lane="6" entrytime="00:01:32.15" entrycourse="SCM" />
                <RESULT eventid="1326" status="DNS" swimtime="00:00:00.00" resultid="2787" heatid="5126" lane="2" />
                <RESULT eventid="10329" status="DNS" swimtime="00:00:00.00" resultid="10446" heatid="10344" lane="4" entrytime="00:00:36.64" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="De Almeida Dias" birthdate="2012-02-18" gender="F" nation="BRA" license="369262" swrid="5588638" athleteid="2323" externalid="369262" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="331" swimtime="00:00:35.23" resultid="2324" heatid="4657" lane="1" />
                <RESULT eventid="1077" points="345" swimtime="00:00:35.99" resultid="2325" heatid="4721" lane="3" entrytime="00:00:35.23" entrycourse="SCM" />
                <RESULT eventid="1165" points="372" swimtime="00:01:16.28" resultid="2326" heatid="4914" lane="2" entrytime="00:01:15.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="478" swimtime="00:02:21.06" resultid="2327" heatid="4895" lane="3" entrytime="00:02:22.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                    <SPLIT distance="100" swimtime="00:01:08.71" />
                    <SPLIT distance="150" swimtime="00:01:45.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="398" swimtime="00:00:31.15" resultid="2328" heatid="5096" lane="5" entrytime="00:00:30.28" entrycourse="SCM" />
                <RESULT eventid="1301" points="336" swimtime="00:00:40.78" resultid="2329" heatid="5037" lane="2" />
                <RESULT eventid="4411" points="304" swimtime="00:00:36.24" resultid="5391" heatid="4680" lane="5" />
                <RESULT eventid="4417" points="351" swimtime="00:00:35.77" resultid="5421" heatid="4731" lane="5" />
                <RESULT eventid="4419" points="329" swimtime="00:00:36.55" resultid="5425" heatid="4742" lane="3" />
                <RESULT eventid="5801" points="323" swimtime="00:00:41.34" resultid="10100" heatid="6068" lane="4" />
                <RESULT eventid="5804" points="399" swimtime="00:00:31.13" resultid="10197" heatid="6054" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Da Cunha Souza" birthdate="2013-09-17" gender="M" nation="BRA" license="376975" swrid="5588618" athleteid="2489" externalid="376975" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="117" swimtime="00:00:44.36" resultid="2490" heatid="4775" lane="1" entrytime="00:00:43.89" entrycourse="SCM" />
                <RESULT eventid="1105" points="129" swimtime="00:00:43.74" resultid="2491" heatid="4828" lane="3" />
                <RESULT eventid="1227" points="187" swimtime="00:02:53.57" resultid="2492" heatid="4966" lane="1" entrytime="00:03:02.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.17" />
                    <SPLIT distance="100" swimtime="00:01:23.97" />
                    <SPLIT distance="150" swimtime="00:02:09.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="180" swimtime="00:01:19.38" resultid="2493" heatid="5004" lane="2" entrytime="00:01:21.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="132" swimtime="00:00:48.88" resultid="2495" heatid="5148" lane="3" entrytime="00:00:54.82" entrycourse="SCM" />
                <RESULT eventid="10332" points="195" swimtime="00:00:34.75" resultid="10424" heatid="10350" lane="4" entrytime="00:00:36.07" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Muxfeldt" birthdate="2011-05-13" gender="F" nation="BRA" license="366903" swrid="5602563" athleteid="2274" externalid="366903" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="266" swimtime="00:00:37.89" resultid="2275" heatid="4661" lane="6" />
                <RESULT eventid="1077" points="317" swimtime="00:00:37.00" resultid="2276" heatid="4712" lane="3" />
                <RESULT eventid="1119" points="326" swimtime="00:02:52.73" resultid="2277" heatid="4874" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.70" />
                    <SPLIT distance="100" swimtime="00:02:09.91" />
                    <SPLIT distance="150" swimtime="00:02:52.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="193" swimtime="00:01:33.50" resultid="2278" heatid="4899" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="385" swimtime="00:00:31.51" resultid="2279" heatid="5093" lane="7" entrytime="00:00:32.53" entrycourse="SCM" />
                <RESULT eventid="1301" points="335" swimtime="00:00:40.83" resultid="2280" heatid="5044" lane="5" entrytime="00:00:42.38" entrycourse="SCM" />
                <RESULT eventid="4417" points="300" swimtime="00:00:37.68" resultid="5431" heatid="4733" lane="6" />
                <RESULT eventid="5801" points="315" swimtime="00:00:41.69" resultid="10158" heatid="6070" lane="5" />
                <RESULT eventid="5804" points="400" swimtime="00:00:31.10" resultid="10198" heatid="6056" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Toscani Kim" birthdate="2015-10-02" gender="F" nation="BRA" license="397276" swrid="5641778" athleteid="2823" externalid="397276" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="201" swimtime="00:00:41.57" resultid="2824" heatid="4650" lane="4" entrytime="00:00:46.83" entrycourse="SCM" />
                <RESULT eventid="1074" points="165" swimtime="00:00:46.00" resultid="2825" heatid="4702" lane="1" entrytime="00:00:46.39" entrycourse="SCM" />
                <RESULT eventid="1129" points="197" swimtime="00:01:47.14" resultid="2826" heatid="4881" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="139" swimtime="00:01:44.27" resultid="2827" heatid="4898" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="192" swimtime="00:00:49.12" resultid="2828" heatid="5025" lane="1" entrytime="00:00:51.49" entrycourse="SCM" />
                <RESULT eventid="1311" points="177" swimtime="00:00:40.80" resultid="2829" heatid="5076" lane="8" entrytime="00:00:40.77" entrycourse="SCM" />
                <RESULT eventid="4409" points="209" swimtime="00:00:41.06" resultid="5365" heatid="4655" lane="3" />
                <RESULT eventid="4415" points="159" swimtime="00:00:46.53" resultid="5398" heatid="4706" lane="3" />
                <RESULT eventid="4433" points="203" swimtime="00:00:48.23" resultid="10080" heatid="5029" lane="2" />
                <RESULT eventid="4439" points="187" swimtime="00:00:40.05" resultid="10179" heatid="6048" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Marie Silva" birthdate="2014-08-24" gender="F" nation="BRA" license="391025" swrid="5602556" athleteid="2697" externalid="391025" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" status="DNS" swimtime="00:00:00.00" resultid="2698" heatid="4649" lane="3" entrytime="00:00:53.26" entrycourse="SCM" />
                <RESULT eventid="1074" status="DNS" swimtime="00:00:00.00" resultid="2699" heatid="4697" lane="5" />
                <RESULT eventid="1129" status="DNS" swimtime="00:00:00.00" resultid="2700" heatid="4882" lane="3" />
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="2701" heatid="4906" lane="6" />
                <RESULT eventid="1298" status="DNS" swimtime="00:00:00.00" resultid="2702" heatid="5024" lane="2" entrytime="00:00:55.80" entrycourse="SCM" />
                <RESULT eventid="1311" status="DNS" swimtime="00:00:00.00" resultid="2703" heatid="5075" lane="6" entrytime="00:00:41.68" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Schiavon" birthdate="2010-05-03" gender="M" nation="BRA" license="356354" swrid="5600256" athleteid="2218" externalid="356354" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="2219" heatid="4772" lane="5" />
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="2220" heatid="4827" lane="5" />
                <RESULT eventid="1227" points="378" swimtime="00:02:17.43" resultid="2221" heatid="4965" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                    <SPLIT distance="100" swimtime="00:01:05.82" />
                    <SPLIT distance="150" swimtime="00:01:43.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="331" swimtime="00:01:04.81" resultid="2222" heatid="5000" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" status="DNS" swimtime="00:00:00.00" resultid="2224" heatid="5147" lane="8" />
                <RESULT eventid="10332" status="DNS" swimtime="00:00:00.00" resultid="10403" heatid="10348" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="De Macedo Martynychen" birthdate="2015-06-12" gender="F" nation="BRA" license="399681" swrid="5652885" athleteid="2837" externalid="399681" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" status="DNS" swimtime="00:00:00.00" resultid="2838" heatid="4648" lane="6" entrytime="00:01:02.44" entrycourse="SCM" />
                <RESULT eventid="1074" status="DNS" swimtime="00:00:00.00" resultid="2839" heatid="4698" lane="2" entrytime="00:00:57.10" entrycourse="SCM" />
                <RESULT eventid="1165" points="65" swimtime="00:02:15.97" resultid="2840" heatid="4904" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1153" points="91" swimtime="00:02:00.11" resultid="2841" heatid="4898" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="89" swimtime="00:01:03.50" resultid="2842" heatid="5020" lane="1" />
                <RESULT eventid="1311" points="87" swimtime="00:00:51.68" resultid="2843" heatid="5071" lane="3" entrytime="00:00:51.80" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Szpak De Vasconcelos" birthdate="2012-06-29" gender="M" nation="BRA" license="369271" swrid="5588928" athleteid="2356" externalid="369271" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="219" swimtime="00:00:36.05" resultid="2357" heatid="4766" lane="4" />
                <RESULT eventid="1105" points="235" swimtime="00:00:35.79" resultid="2358" heatid="4839" lane="5" entrytime="00:00:36.02" entrycourse="SCM" />
                <RESULT eventid="1213" points="299" swimtime="00:01:22.62" resultid="2359" heatid="4953" lane="2" entrytime="00:01:23.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="234" swimtime="00:01:18.32" resultid="2360" heatid="4979" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="282" swimtime="00:00:38.02" resultid="2362" heatid="5154" lane="3" entrytime="00:00:38.19" entrycourse="SCM" />
                <RESULT eventid="4429" points="247" swimtime="00:00:35.21" resultid="5522" heatid="4854" lane="3" />
                <RESULT eventid="4431" points="244" swimtime="00:00:35.38" resultid="5528" heatid="4865" lane="3" />
                <RESULT eventid="5807" points="297" swimtime="00:00:37.39" resultid="10276" heatid="6038" lane="5" />
                <RESULT eventid="10332" points="316" swimtime="00:00:29.59" resultid="10416" heatid="10356" lane="8" entrytime="00:00:29.92" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Rampazzo" birthdate="2013-02-18" gender="M" nation="BRA" license="400269" swrid="5748679" athleteid="3033" externalid="400269" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="164" swimtime="00:00:39.71" resultid="3034" heatid="4773" lane="3" />
                <RESULT eventid="1105" points="169" swimtime="00:00:39.97" resultid="3035" heatid="4826" lane="4" />
                <RESULT eventid="1213" points="268" swimtime="00:01:25.72" resultid="3036" heatid="4952" lane="4" entrytime="00:01:34.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="232" swimtime="00:03:15.49" resultid="3037" heatid="4993" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.62" />
                    <SPLIT distance="100" swimtime="00:01:33.41" />
                    <SPLIT distance="150" swimtime="00:02:26.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="270" swimtime="00:00:38.56" resultid="3039" heatid="5152" lane="2" entrytime="00:00:41.38" entrycourse="SCM" />
                <RESULT eventid="5807" points="272" swimtime="00:00:38.48" resultid="10269" heatid="6036" lane="4" />
                <RESULT eventid="10332" points="263" swimtime="00:00:31.44" resultid="10463" heatid="10352" lane="4" entrytime="00:00:33.65" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Steven" lastname="Matheussi Viana E Silva" birthdate="2012-05-03" gender="M" nation="BRA" license="376986" swrid="5588810" athleteid="2552" externalid="376986" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="229" swimtime="00:00:35.52" resultid="2553" heatid="4777" lane="4" entrytime="00:00:36.79" entrycourse="SCM" />
                <RESULT eventid="1105" points="154" swimtime="00:00:41.17" resultid="2554" heatid="4829" lane="5" />
                <RESULT eventid="1213" points="263" swimtime="00:01:26.20" resultid="2555" heatid="4953" lane="6" entrytime="00:01:29.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="263" swimtime="00:03:07.53" resultid="2556" heatid="4993" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.42" />
                    <SPLIT distance="100" swimtime="00:01:29.16" />
                    <SPLIT distance="150" swimtime="00:02:17.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="271" swimtime="00:00:38.55" resultid="2558" heatid="5152" lane="7" entrytime="00:00:39.87" entrycourse="SCM" />
                <RESULT eventid="5807" points="267" swimtime="00:00:38.70" resultid="10274" heatid="6038" lane="3" />
                <RESULT eventid="10332" points="275" swimtime="00:00:30.98" resultid="10430" heatid="10352" lane="6" entrytime="00:00:34.84" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Bau Santos" birthdate="2015-05-28" gender="M" nation="BRA" license="417451" athleteid="3066" externalid="417451" level="CLBO">
              <RESULTS>
                <RESULT eventid="1102" status="DNS" swimtime="00:00:00.00" resultid="3067" heatid="4811" lane="6" />
                <RESULT eventid="1213" status="DNS" swimtime="00:00:00.00" resultid="3068" heatid="4947" lane="1" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="3069" heatid="4999" lane="5" />
                <RESULT eventid="1326" status="DNS" swimtime="00:00:00.00" resultid="3071" heatid="5124" lane="3" />
                <RESULT eventid="10329" status="DNS" swimtime="00:00:00.00" resultid="10467" heatid="10341" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Azevedo Alanis" birthdate="2013-12-07" gender="M" nation="BRA" license="376991" swrid="5588540" athleteid="2531" externalid="376991" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="109" swimtime="00:00:45.44" resultid="2532" heatid="4772" lane="4" />
                <RESULT eventid="1105" points="123" swimtime="00:00:44.40" resultid="2533" heatid="4833" lane="4" />
                <RESULT eventid="1213" points="147" swimtime="00:01:44.58" resultid="2534" heatid="4952" lane="6" entrytime="00:01:43.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1263" points="151" swimtime="00:03:45.44" resultid="2535" heatid="4993" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.32" />
                    <SPLIT distance="100" swimtime="00:01:49.62" />
                    <SPLIT distance="150" swimtime="00:02:47.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="145" swimtime="00:00:47.42" resultid="2537" heatid="5151" lane="7" entrytime="00:00:48.80" entrycourse="SCM" />
                <RESULT eventid="10332" points="152" swimtime="00:00:37.70" resultid="10428" heatid="10350" lane="7" entrytime="00:00:39.31" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martina" lastname="Mayer Paludetto" birthdate="2012-10-30" gender="F" nation="BRA" license="369264" swrid="5588811" athleteid="2330" externalid="369264" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="386" swimtime="00:00:33.46" resultid="2331" heatid="4670" lane="3" entrytime="00:00:35.81" entrycourse="SCM" />
                <RESULT eventid="1077" points="373" swimtime="00:00:35.05" resultid="2332" heatid="4721" lane="1" entrytime="00:00:36.82" entrycourse="SCM" />
                <RESULT eventid="1165" points="395" swimtime="00:01:14.81" resultid="2333" heatid="4913" lane="3" entrytime="00:01:20.98" entrycourse="SCM" />
                <RESULT eventid="1143" points="496" swimtime="00:02:19.34" resultid="2334" heatid="4893" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="417" swimtime="00:00:30.67" resultid="2335" heatid="5096" lane="3" entrytime="00:00:29.80" entrycourse="SCM" />
                <RESULT eventid="1301" points="341" swimtime="00:00:40.57" resultid="2336" heatid="5042" lane="6" entrytime="00:00:44.08" entrycourse="SCM" />
                <RESULT eventid="4411" points="379" swimtime="00:00:33.67" resultid="5389" heatid="4680" lane="3" />
                <RESULT eventid="4413" points="354" swimtime="00:00:34.45" resultid="5395" heatid="4691" lane="3" />
                <RESULT eventid="4417" points="390" swimtime="00:00:34.54" resultid="5418" heatid="4731" lane="2" />
                <RESULT eventid="4419" points="367" swimtime="00:00:35.26" resultid="5424" heatid="4742" lane="2" />
                <RESULT eventid="5801" points="336" swimtime="00:00:40.80" resultid="10099" heatid="6068" lane="3" />
                <RESULT eventid="5804" points="439" swimtime="00:00:30.16" resultid="10196" heatid="6054" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Zagonel Krempel" birthdate="2015-07-27" gender="F" nation="BRA" license="406962" swrid="5717305" athleteid="2977" externalid="406962" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" status="DNS" swimtime="00:00:00.00" resultid="2978" heatid="4646" lane="5" />
                <RESULT eventid="1074" status="DNS" swimtime="00:00:00.00" resultid="2979" heatid="4698" lane="4" entrytime="00:00:57.09" entrycourse="SCM" />
                <RESULT eventid="1129" status="DNS" swimtime="00:00:00.00" resultid="2980" heatid="4882" lane="5" />
                <RESULT eventid="1189" status="DNS" swimtime="00:00:00.00" resultid="2981" heatid="4926" lane="2" entrytime="00:02:03.97" entrycourse="SCM" />
                <RESULT eventid="1298" status="DNS" swimtime="00:00:00.00" resultid="2982" heatid="5021" lane="5" entrytime="00:01:09.08" entrycourse="SCM" />
                <RESULT eventid="1311" status="DNS" swimtime="00:00:00.00" resultid="2983" heatid="5071" lane="4" entrytime="00:00:51.96" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Mattioli" birthdate="2011-10-22" gender="F" nation="BRA" license="366896" swrid="5602559" athleteid="2253" externalid="366896" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="316" swimtime="00:00:35.79" resultid="2254" heatid="4659" lane="1" />
                <RESULT eventid="1077" points="321" swimtime="00:00:36.86" resultid="2255" heatid="4712" lane="2" />
                <RESULT eventid="1129" points="439" swimtime="00:01:22.03" resultid="2256" heatid="4886" lane="1" entrytime="00:01:31.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="441" swimtime="00:02:56.69" resultid="2257" heatid="4922" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.77" />
                    <SPLIT distance="100" swimtime="00:01:24.89" />
                    <SPLIT distance="150" swimtime="00:02:11.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="374" swimtime="00:00:31.82" resultid="2258" heatid="5094" lane="5" entrytime="00:00:31.18" entrycourse="SCM" />
                <RESULT eventid="1301" points="416" swimtime="00:00:37.99" resultid="2259" heatid="5036" lane="7" />
                <RESULT eventid="4417" points="351" swimtime="00:00:35.77" resultid="5429" heatid="4733" lane="4" />
                <RESULT eventid="5801" points="393" swimtime="00:00:38.72" resultid="10154" heatid="6070" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcela" lastname="Tallao Benke" birthdate="2014-10-07" gender="F" nation="BRA" license="382075" swrid="5602586" athleteid="2566" externalid="382075" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="292" swimtime="00:00:36.73" resultid="2567" heatid="4651" lane="3" entrytime="00:00:39.27" entrycourse="SCM" />
                <RESULT eventid="1074" points="242" swimtime="00:00:40.50" resultid="2568" heatid="4696" lane="5" />
                <RESULT eventid="1129" points="246" swimtime="00:01:39.49" resultid="2569" heatid="4882" lane="6" />
                <RESULT eventid="1153" points="241" swimtime="00:01:26.76" resultid="2570" heatid="4899" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="251" swimtime="00:00:44.93" resultid="2571" heatid="5025" lane="4" entrytime="00:00:45.52" entrycourse="SCM" />
                <RESULT eventid="1311" points="296" swimtime="00:00:34.40" resultid="2572" heatid="5076" lane="4" entrytime="00:00:34.87" entrycourse="SCM" />
                <RESULT eventid="4409" points="294" swimtime="00:00:36.64" resultid="5371" heatid="4656" lane="1" />
                <RESULT eventid="4415" points="255" swimtime="00:00:39.80" resultid="5402" heatid="4707" lane="1" />
                <RESULT eventid="4433" points="256" swimtime="00:00:44.65" resultid="10086" heatid="6064" lane="2" />
                <RESULT eventid="4439" points="296" swimtime="00:00:34.38" resultid="10182" heatid="6050" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio" lastname="Carcereri Navarro" birthdate="2013-12-19" gender="M" nation="BRA" license="376962" swrid="5588576" athleteid="2475" externalid="376962" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="175" swimtime="00:00:38.83" resultid="2476" heatid="4776" lane="1" entrytime="00:00:40.01" entrycourse="SCM" />
                <RESULT eventid="1105" points="116" swimtime="00:00:45.31" resultid="2477" heatid="4829" lane="1" />
                <RESULT comment="SW 7.4 - Movimentos das pernas não simultâneos., SW 7.5 - Pé esquerdo não virado para fora durante a parte propulsora da pernada (fim do ciclo)." eventid="1213" status="DSQ" swimtime="00:01:38.67" resultid="2478" heatid="4952" lane="1" entrytime="00:01:42.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1237" points="137" swimtime="00:01:32.64" resultid="2479" heatid="4972" lane="6" entrytime="00:01:37.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="157" swimtime="00:00:46.21" resultid="2481" heatid="5151" lane="3" entrytime="00:00:44.44" entrycourse="SCM" />
                <RESULT eventid="10332" points="195" swimtime="00:00:34.72" resultid="10423" heatid="10351" lane="7" entrytime="00:00:36.63" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Schmidt Wozniaki" birthdate="2012-07-07" gender="M" nation="BRA" license="376963" swrid="5588905" athleteid="5256" externalid="376963" level="CLBO">
              <RESULTS>
                <RESULT eventid="1329" points="158" swimtime="00:00:46.07" resultid="5258" heatid="5139" lane="1" />
                <RESULT eventid="1092" points="131" swimtime="00:00:42.78" resultid="5259" heatid="4762" lane="5" />
                <RESULT eventid="1105" points="113" swimtime="00:00:45.68" resultid="5260" heatid="5253" lane="5" />
                <RESULT eventid="10332" points="197" swimtime="00:00:34.64" resultid="10542" heatid="10347" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Fernandes" birthdate="2010-03-13" gender="M" nation="BRA" license="339266" swrid="5588695" athleteid="2608" externalid="339266" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="403" swimtime="00:00:29.43" resultid="2609" heatid="4774" lane="5" />
                <RESULT eventid="1105" points="348" swimtime="00:00:31.41" resultid="2610" heatid="4841" lane="2" entrytime="00:00:30.36" entrycourse="SCM" />
                <RESULT eventid="1227" points="499" swimtime="00:02:05.25" resultid="2611" heatid="4963" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                    <SPLIT distance="100" swimtime="00:01:01.47" />
                    <SPLIT distance="150" swimtime="00:01:33.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="504" swimtime="00:00:56.33" resultid="2612" heatid="5010" lane="2" entrytime="00:00:58.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="354" swimtime="00:00:35.24" resultid="2614" heatid="5138" lane="3" />
                <RESULT eventid="4423" points="392" swimtime="00:00:29.70" resultid="5538" heatid="4798" lane="1" />
                <RESULT eventid="4425" points="377" swimtime="00:00:30.10" resultid="5544" heatid="4807" lane="1" />
                <RESULT eventid="4429" points="335" swimtime="00:00:31.83" resultid="5576" heatid="4858" lane="1" />
                <RESULT eventid="4431" points="380" swimtime="00:00:30.51" resultid="5582" heatid="4867" lane="1" />
                <RESULT eventid="5807" points="286" swimtime="00:00:37.83" resultid="10289" heatid="6042" lane="5" />
                <RESULT eventid="10332" points="476" swimtime="00:00:25.81" resultid="10435" heatid="10360" lane="7" entrytime="00:00:26.41" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Fernandes  Dos Reis" birthdate="2012-09-18" gender="M" nation="BRA" license="369279" swrid="5588696" athleteid="2398" externalid="369279" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="255" swimtime="00:00:34.29" resultid="2399" heatid="4778" lane="4" entrytime="00:00:33.82" entrycourse="SCM" />
                <RESULT eventid="1105" points="174" swimtime="00:00:39.60" resultid="2400" heatid="4836" lane="3" entrytime="00:00:39.91" entrycourse="SCM" />
                <RESULT eventid="1237" points="235" swimtime="00:01:17.35" resultid="2401" heatid="4973" lane="1" entrytime="00:01:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="254" swimtime="00:01:10.75" resultid="2402" heatid="5007" lane="1" entrytime="00:01:08.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente., Na volta dos 25m." eventid="1329" status="DSQ" swimtime="00:00:47.53" resultid="2404" heatid="5150" lane="3" entrytime="00:00:45.93" entrycourse="SCM" />
                <RESULT eventid="4423" points="249" swimtime="00:00:34.55" resultid="5498" heatid="4794" lane="6" />
                <RESULT eventid="4425" points="249" swimtime="00:00:34.55" resultid="9034" heatid="9999" lane="3" />
                <RESULT eventid="10332" points="256" swimtime="00:00:31.72" resultid="10419" heatid="10353" lane="3" entrytime="00:00:31.99" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Vanzo Assumpcao" birthdate="2012-05-15" gender="M" nation="BRA" license="369258" swrid="5588942" athleteid="2309" externalid="369258" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="360" swimtime="00:00:30.55" resultid="2310" heatid="4779" lane="6" entrytime="00:00:32.82" entrycourse="SCM" />
                <RESULT eventid="1105" points="275" swimtime="00:00:33.96" resultid="2311" heatid="4840" lane="1" entrytime="00:00:34.28" entrycourse="SCM" />
                <RESULT eventid="1203" points="316" swimtime="00:02:34.99" resultid="2312" heatid="4943" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                    <SPLIT distance="100" swimtime="00:01:17.43" />
                    <SPLIT distance="150" swimtime="00:01:56.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1227" points="368" swimtime="00:02:18.65" resultid="2313" heatid="4967" lane="6" entrytime="00:02:35.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.80" />
                    <SPLIT distance="100" swimtime="00:01:08.31" />
                    <SPLIT distance="150" swimtime="00:01:43.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="222" swimtime="00:00:41.20" resultid="2315" heatid="5138" lane="4" />
                <RESULT eventid="4423" points="364" swimtime="00:00:30.44" resultid="5493" heatid="4794" lane="1" />
                <RESULT eventid="4429" points="285" swimtime="00:00:33.56" resultid="5520" heatid="4854" lane="1" />
                <RESULT eventid="4431" points="283" swimtime="00:00:33.65" resultid="5526" heatid="4865" lane="1" />
                <RESULT eventid="4425" points="322" swimtime="00:00:31.70" resultid="5603" heatid="4805" lane="1" />
                <RESULT eventid="5807" points="207" swimtime="00:00:42.14" resultid="10278" heatid="6038" lane="7" />
                <RESULT eventid="10332" points="355" swimtime="00:00:28.45" resultid="10411" heatid="10354" lane="4" entrytime="00:00:31.64" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Fontana" birthdate="2011-12-29" gender="M" nation="BRA" license="366897" swrid="5602539" athleteid="2260" externalid="366897" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="170" swimtime="00:00:39.26" resultid="2261" heatid="4765" lane="1" />
                <RESULT eventid="1105" points="157" swimtime="00:00:40.94" resultid="2262" heatid="4827" lane="3" />
                <RESULT eventid="1213" points="187" swimtime="00:01:36.56" resultid="2263" heatid="4952" lane="2" entrytime="00:01:36.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="153" swimtime="00:01:30.29" resultid="2264" heatid="4984" lane="3" entrytime="00:01:28.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="204" swimtime="00:00:42.36" resultid="2266" heatid="5143" lane="2" />
                <RESULT eventid="10332" points="212" swimtime="00:00:33.77" resultid="10408" heatid="10351" lane="6" entrytime="00:00:35.71" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Cabrera Cirino Dos Santos" birthdate="2013-03-30" gender="M" nation="BRA" license="376990" swrid="5588570" athleteid="2538" externalid="376990" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="173" swimtime="00:00:39.03" resultid="2539" heatid="4775" lane="6" entrytime="00:00:46.02" entrycourse="SCM" />
                <RESULT eventid="1105" points="160" swimtime="00:00:40.71" resultid="2540" heatid="4835" lane="4" entrytime="00:00:44.67" entrycourse="SCM" />
                <RESULT eventid="1227" points="238" swimtime="00:02:40.29" resultid="2541" heatid="4966" lane="5" entrytime="00:02:54.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                    <SPLIT distance="100" swimtime="00:01:18.59" />
                    <SPLIT distance="150" swimtime="00:01:59.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="207" swimtime="00:01:15.71" resultid="2542" heatid="5005" lane="5" entrytime="00:01:15.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" status="DNS" swimtime="00:00:00.00" resultid="2544" heatid="5147" lane="2" />
                <RESULT eventid="4429" points="183" swimtime="00:00:38.89" resultid="5515" heatid="4852" lane="5" />
                <RESULT eventid="10332" points="211" swimtime="00:00:33.82" resultid="10429" heatid="10352" lane="2" entrytime="00:00:34.29" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olavo" lastname="Valduga Artigas" birthdate="2012-06-26" gender="M" nation="BRA" license="369270" swrid="5588941" athleteid="2351" externalid="369270" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="113" swimtime="00:00:44.94" resultid="2352" heatid="4766" lane="3" />
                <RESULT eventid="1105" points="106" swimtime="00:00:46.66" resultid="2353" heatid="4827" lane="6" />
                <RESULT eventid="1329" points="143" swimtime="00:00:47.63" resultid="2355" heatid="5151" lane="5" entrytime="00:00:45.16" entrycourse="SCM" />
                <RESULT eventid="10332" points="179" swimtime="00:00:35.77" resultid="10415" heatid="10350" lane="5" entrytime="00:00:36.31" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Guimaraes Mesquita" birthdate="2015-10-05" gender="F" nation="BRA" license="393263" swrid="5616444" athleteid="2774" externalid="393263" level="CLBO">
              <RESULTS>
                <RESULT comment="SW 8.3 - Movimento de pernada de peito.&#10;&#10;&#10;&#10;&#10;&#10;&#10;" eventid="1061" status="DSQ" swimtime="00:01:20.86" resultid="2775" heatid="4647" lane="6" entrytime="00:01:35.32" entrycourse="SCM" />
                <RESULT eventid="1074" points="66" swimtime="00:01:02.34" resultid="2776" heatid="4697" lane="4" entrytime="00:01:05.64" entrycourse="SCM" />
                <RESULT eventid="1129" points="78" swimtime="00:02:25.73" resultid="2777" heatid="4883" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="65" swimtime="00:02:16.50" resultid="2778" heatid="4910" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="72" swimtime="00:01:07.89" resultid="2779" heatid="5021" lane="1" entrytime="00:01:10.43" entrycourse="SCM" />
                <RESULT eventid="1311" points="60" swimtime="00:00:58.32" resultid="2780" heatid="5071" lane="6" entrytime="00:01:00.49" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Cecilia Carvalho" birthdate="2014-10-30" gender="F" nation="BRA" license="391021" swrid="5602525" athleteid="2676" externalid="391021" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" points="134" swimtime="00:00:47.61" resultid="2677" heatid="4650" lane="5" entrytime="00:00:49.98" entrycourse="SCM" />
                <RESULT eventid="1074" points="138" swimtime="00:00:48.82" resultid="2678" heatid="4700" lane="4" entrytime="00:00:50.79" entrycourse="SCM" />
                <RESULT eventid="1129" points="99" swimtime="00:02:14.67" resultid="2679" heatid="4883" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="110" swimtime="00:01:54.36" resultid="2680" heatid="4910" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="98" swimtime="00:01:01.40" resultid="2681" heatid="5021" lane="3" entrytime="00:01:06.32" entrycourse="SCM" />
                <RESULT eventid="1311" points="215" swimtime="00:00:38.24" resultid="2682" heatid="5076" lane="7" entrytime="00:00:41.24" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Fontolan Gomes" birthdate="2010-07-02" gender="M" nation="BRA" license="356245" swrid="5588705" athleteid="2204" externalid="356245" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="193" swimtime="00:00:37.63" resultid="2205" heatid="4765" lane="4" />
                <RESULT eventid="1105" points="259" swimtime="00:00:34.65" resultid="2206" heatid="4840" lane="6" entrytime="00:00:34.55" entrycourse="SCM" />
                <RESULT eventid="1213" points="222" swimtime="00:01:31.25" resultid="2207" heatid="4952" lane="3" entrytime="00:01:32.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="324" swimtime="00:01:10.31" resultid="2208" heatid="4986" lane="1" entrytime="00:01:10.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="209" swimtime="00:00:41.98" resultid="2210" heatid="5146" lane="1" />
                <RESULT eventid="4429" points="266" swimtime="00:00:34.36" resultid="5579" heatid="4858" lane="4" />
                <RESULT eventid="10332" points="300" swimtime="00:00:30.10" resultid="10401" heatid="10348" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alan" lastname="Batista Grise" birthdate="2014-03-27" gender="M" nation="BRA" license="391007" swrid="5602513" athleteid="2622" externalid="391007" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" status="DNS" swimtime="00:00:00.00" resultid="2623" heatid="4751" lane="1" />
                <RESULT eventid="1102" status="DNS" swimtime="00:00:00.00" resultid="2624" heatid="4810" lane="2" />
                <RESULT eventid="1249" status="DNS" swimtime="00:00:00.00" resultid="2625" heatid="4979" lane="1" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="2626" heatid="5001" lane="4" entrytime="00:01:50.70" entrycourse="SCM" />
                <RESULT eventid="1326" status="DNS" swimtime="00:00:00.00" resultid="2628" heatid="5128" lane="5" entrytime="00:01:02.87" entrycourse="SCM" />
                <RESULT eventid="10329" status="DNS" swimtime="00:00:00.00" resultid="10436" heatid="10342" lane="5" entrytime="00:00:46.96" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="De Moraes" birthdate="2014-09-18" gender="M" nation="BRA" license="391024" swrid="5602529" athleteid="2690" externalid="391024" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="185" swimtime="00:00:38.17" resultid="2691" heatid="4756" lane="2" entrytime="00:00:40.46" entrycourse="SCM" />
                <RESULT eventid="1102" points="163" swimtime="00:00:40.42" resultid="2692" heatid="4817" lane="5" entrytime="00:00:41.49" entrycourse="SCM" />
                <RESULT eventid="1213" points="154" swimtime="00:01:43.09" resultid="2693" heatid="4947" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="159" swimtime="00:01:29.16" resultid="2694" heatid="4979" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="162" swimtime="00:00:45.74" resultid="2696" heatid="5131" lane="5" entrytime="00:00:50.20" entrycourse="SCM" />
                <RESULT eventid="4421" points="185" swimtime="00:00:38.12" resultid="5469" heatid="4761" lane="1" />
                <RESULT eventid="4427" points="171" swimtime="00:00:39.80" resultid="5506" heatid="4822" lane="2" />
                <RESULT eventid="4445" points="172" swimtime="00:00:44.80" resultid="10315" heatid="6034" lane="5" />
                <RESULT eventid="10329" points="256" swimtime="00:00:31.74" resultid="10442" heatid="10345" lane="3" entrytime="00:00:32.45" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Hadad" birthdate="2015-09-09" gender="M" nation="BRA" license="406740" swrid="5717272" athleteid="2886" externalid="406740" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" status="DNS" swimtime="00:00:00.00" resultid="2887" heatid="4750" lane="1" />
                <RESULT eventid="1102" points="74" swimtime="00:00:52.58" resultid="2888" heatid="4813" lane="4" entrytime="00:00:57.64" entrycourse="SCM" />
                <RESULT eventid="1249" points="60" swimtime="00:02:02.84" resultid="2889" heatid="4982" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1237" points="49" swimtime="00:02:10.12" resultid="2890" heatid="4970" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="57" swimtime="00:01:04.78" resultid="2892" heatid="5127" lane="3" entrytime="00:01:08.06" entrycourse="SCM" />
                <RESULT eventid="10329" points="99" swimtime="00:00:43.50" resultid="10451" heatid="10342" lane="1" entrytime="00:00:47.28" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Saporiti Salvi" birthdate="2013-06-28" gender="M" nation="BRA" license="377032" swrid="5588896" athleteid="2517" externalid="377032" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="173" swimtime="00:00:38.96" resultid="2518" heatid="4776" lane="2" entrytime="00:00:38.27" entrycourse="SCM" />
                <RESULT eventid="1105" points="159" swimtime="00:00:40.75" resultid="2519" heatid="4825" lane="3" />
                <RESULT eventid="1237" points="170" swimtime="00:01:26.15" resultid="2520" heatid="4972" lane="5" entrytime="00:01:27.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="218" swimtime="00:01:14.43" resultid="2521" heatid="5005" lane="2" entrytime="00:01:15.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="143" swimtime="00:00:47.71" resultid="2523" heatid="5148" lane="8" entrytime="00:00:49.56" entrycourse="SCM" />
                <RESULT eventid="10332" points="226" swimtime="00:00:33.05" resultid="10426" heatid="10351" lane="3" entrytime="00:00:35.17" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Shwetz Clivatti" birthdate="2015-03-05" gender="M" nation="BRA" license="406963" swrid="5717297" athleteid="2984" externalid="406963" level="CLBO">
              <RESULTS>
                <RESULT eventid="1102" status="DNS" swimtime="00:00:00.00" resultid="2985" heatid="4812" lane="5" entrytime="00:01:07.34" entrycourse="SCM" />
                <RESULT eventid="1213" status="DNS" swimtime="00:00:00.00" resultid="2986" heatid="4947" lane="3" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="2987" heatid="5001" lane="2" entrytime="00:02:10.13" entrycourse="SCM" />
                <RESULT eventid="1326" status="DNS" swimtime="00:00:00.00" resultid="2989" heatid="5127" lane="5" entrytime="00:01:15.50" entrycourse="SCM" />
                <RESULT eventid="10329" status="DNS" swimtime="00:00:00.00" resultid="10459" heatid="10340" lane="5" entrytime="00:01:01.73" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Xavier Jardim" birthdate="2012-01-23" gender="M" nation="BRA" license="369259" swrid="5641781" athleteid="2316" externalid="369259" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="240" swimtime="00:00:34.99" resultid="2317" heatid="4776" lane="5" entrytime="00:00:39.40" entrycourse="SCM" />
                <RESULT eventid="1105" points="184" swimtime="00:00:38.85" resultid="2318" heatid="4837" lane="2" entrytime="00:00:38.73" entrycourse="SCM" />
                <RESULT eventid="1237" points="171" swimtime="00:01:25.96" resultid="2319" heatid="4972" lane="2" entrytime="00:01:26.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="259" swimtime="00:01:10.26" resultid="2320" heatid="5007" lane="6" entrytime="00:01:08.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" status="DNS" swimtime="00:00:00.00" resultid="2322" heatid="5146" lane="4" />
                <RESULT eventid="4423" points="237" swimtime="00:00:35.12" resultid="5496" heatid="4794" lane="4" />
                <RESULT eventid="10332" status="DNS" swimtime="00:00:00.00" resultid="10412" heatid="10355" lane="2" entrytime="00:00:31.02" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Alice Silva Gomes Xavier" birthdate="2013-02-25" gender="F" nation="BRA" license="371040" swrid="5717241" athleteid="2963" externalid="371040" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="359" swimtime="00:00:34.30" resultid="2964" heatid="4668" lane="3" entrytime="00:00:39.17" entrycourse="SCM" />
                <RESULT eventid="1077" points="225" swimtime="00:00:41.50" resultid="2965" heatid="4709" lane="1" />
                <RESULT eventid="1129" points="296" swimtime="00:01:33.52" resultid="2966" heatid="4885" lane="3" entrytime="00:01:34.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="272" swimtime="00:03:27.66" resultid="2967" heatid="4920" lane="5" />
                <RESULT eventid="1314" points="351" swimtime="00:00:32.48" resultid="2968" heatid="5093" lane="5" entrytime="00:00:32.12" entrycourse="SCM" />
                <RESULT eventid="1301" points="322" swimtime="00:00:41.36" resultid="2969" heatid="5044" lane="1" entrytime="00:00:41.98" entrycourse="SCM" />
                <RESULT eventid="4413" points="254" swimtime="00:00:38.46" resultid="5375" heatid="4690" lane="1" />
                <RESULT eventid="4411" points="343" swimtime="00:00:34.81" resultid="5381" heatid="4678" lane="1" />
                <RESULT eventid="5801" points="316" swimtime="00:00:41.61" resultid="10091" heatid="6066" lane="1" />
                <RESULT eventid="5804" points="370" swimtime="00:00:31.94" resultid="10190" heatid="6052" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniela" lastname="Alzamora Calado" birthdate="2013-04-26" gender="F" nation="BRA" license="376960" swrid="5588522" athleteid="2461" externalid="376960" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="289" swimtime="00:00:36.85" resultid="2462" heatid="4667" lane="3" entrytime="00:00:40.52" entrycourse="SCM" />
                <RESULT eventid="1077" points="251" swimtime="00:00:39.99" resultid="2463" heatid="4710" lane="6" />
                <RESULT eventid="1179" points="295" swimtime="00:03:22.07" resultid="2464" heatid="4920" lane="4" />
                <RESULT eventid="1189" points="355" swimtime="00:01:10.91" resultid="2465" heatid="4929" lane="6" entrytime="00:01:21.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="392" swimtime="00:00:31.31" resultid="2466" heatid="5092" lane="4" entrytime="00:00:32.63" entrycourse="SCM" />
                <RESULT eventid="1301" points="320" swimtime="00:00:41.47" resultid="2467" heatid="5042" lane="1" entrytime="00:00:43.85" entrycourse="SCM" />
                <RESULT eventid="4411" points="278" swimtime="00:00:37.34" resultid="5384" heatid="4678" lane="4" />
                <RESULT eventid="5801" points="311" swimtime="00:00:41.86" resultid="10093" heatid="6066" lane="3" />
                <RESULT eventid="5804" points="402" swimtime="00:00:31.05" resultid="10186" heatid="6052" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Felipe Canalli" birthdate="2015-12-23" gender="M" nation="BRA" license="406749" swrid="5717261" athleteid="2928" externalid="406749" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="74" swimtime="00:00:51.80" resultid="2929" heatid="4753" lane="3" entrytime="00:01:03.16" entrycourse="SCM" />
                <RESULT eventid="1102" points="56" swimtime="00:00:57.75" resultid="2930" heatid="4812" lane="2" entrytime="00:01:05.26" entrycourse="SCM" />
                <RESULT eventid="1213" points="150" swimtime="00:01:43.95" resultid="2931" heatid="4950" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1237" status="DNS" swimtime="00:00:00.00" resultid="2932" heatid="4969" lane="4" />
                <RESULT eventid="1326" points="150" swimtime="00:00:46.95" resultid="2934" heatid="5130" lane="6" entrytime="00:00:55.35" entrycourse="SCM" />
                <RESULT eventid="4445" points="152" swimtime="00:00:46.69" resultid="10309" heatid="6032" lane="5" />
                <RESULT eventid="10329" points="93" swimtime="00:00:44.41" resultid="10455" heatid="10341" lane="3" entrytime="00:00:51.71" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Galvao" birthdate="2011-03-11" gender="M" nation="BRA" license="381989" swrid="5602541" athleteid="2559" externalid="381989" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="2560" heatid="4769" lane="1" />
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="2561" heatid="4825" lane="4" />
                <RESULT eventid="1237" status="DNS" swimtime="00:00:00.00" resultid="2562" heatid="4970" lane="5" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="2563" heatid="5006" lane="3" entrytime="00:01:09.39" entrycourse="SCM" />
                <RESULT eventid="1329" status="DNS" swimtime="00:00:00.00" resultid="2565" heatid="5144" lane="8" />
                <RESULT eventid="10332" status="DNS" swimtime="00:00:00.00" resultid="10431" heatid="10355" lane="5" entrytime="00:00:31.14" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Miranda Carvalho" birthdate="2015-07-07" gender="F" nation="BRA" license="410200" swrid="5740015" athleteid="3004" externalid="410200" level="CLBO">
              <RESULTS>
                <RESULT eventid="1061" status="DNS" swimtime="00:00:00.00" resultid="3005" heatid="4646" lane="6" />
                <RESULT eventid="1074" status="DNS" swimtime="00:00:00.00" resultid="3006" heatid="4696" lane="4" />
                <RESULT eventid="1165" status="DNS" swimtime="00:00:00.00" resultid="3007" heatid="4907" lane="3" />
                <RESULT eventid="1189" status="DNS" swimtime="00:00:00.00" resultid="3008" heatid="4924" lane="3" />
                <RESULT eventid="1298" status="DNS" swimtime="00:00:00.00" resultid="3009" heatid="5020" lane="5" />
                <RESULT eventid="1311" status="DNS" swimtime="00:00:00.00" resultid="3010" heatid="5072" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gael" lastname="Gluck" birthdate="2011-01-28" gender="M" nation="BRA" license="366891" swrid="5588726" athleteid="2246" externalid="366891" level="CLBO">
              <RESULTS>
                <RESULT eventid="1092" points="342" swimtime="00:00:31.10" resultid="2247" heatid="4765" lane="2" />
                <RESULT eventid="1105" points="218" swimtime="00:00:36.70" resultid="2248" heatid="5253" lane="4" />
                <RESULT eventid="1213" points="390" swimtime="00:01:15.64" resultid="2249" heatid="4953" lane="3" entrytime="00:01:19.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="395" swimtime="00:01:01.11" resultid="2250" heatid="5008" lane="5" entrytime="00:01:04.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1329" points="348" swimtime="00:00:35.47" resultid="2252" heatid="5154" lane="4" entrytime="00:00:36.77" entrycourse="SCM" />
                <RESULT eventid="4423" points="347" swimtime="00:00:30.94" resultid="5533" heatid="4796" lane="5" />
                <RESULT eventid="5807" points="339" swimtime="00:00:35.78" resultid="10281" heatid="6040" lane="4" />
                <RESULT eventid="10332" points="355" swimtime="00:00:28.46" resultid="10407" heatid="10355" lane="7" entrytime="00:00:30.19" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Wolff Contin" birthdate="2015-10-10" gender="M" nation="BRA" license="406745" swrid="5717303" athleteid="2907" externalid="406745" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" status="DNS" swimtime="00:00:00.00" resultid="2908" heatid="4752" lane="3" entrytime="00:01:33.37" entrycourse="SCM" />
                <RESULT eventid="1102" status="DNS" swimtime="00:00:00.00" resultid="2909" heatid="4813" lane="1" entrytime="00:01:03.08" entrycourse="SCM" />
                <RESULT eventid="1249" status="DNS" swimtime="00:00:00.00" resultid="2910" heatid="4981" lane="1" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="2911" heatid="4996" lane="1" />
                <RESULT eventid="1326" status="DNS" swimtime="00:00:00.00" resultid="2913" heatid="5127" lane="1" entrytime="00:01:15.58" entrycourse="SCM" />
                <RESULT eventid="10329" status="DNS" swimtime="00:00:00.00" resultid="10453" heatid="10342" lane="8" entrytime="00:00:51.33" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luisa" lastname="Della Villa Yang" birthdate="2012-10-08" gender="F" nation="BRA" license="369276" swrid="5588653" athleteid="2377" externalid="369276" level="CLBO">
              <RESULTS>
                <RESULT eventid="1064" points="330" swimtime="00:00:35.28" resultid="2378" heatid="4670" lane="4" entrytime="00:00:36.15" entrycourse="SCM" />
                <RESULT eventid="1077" points="276" swimtime="00:00:38.75" resultid="2379" heatid="4718" lane="2" entrytime="00:00:40.39" entrycourse="SCM" />
                <RESULT eventid="1129" points="288" swimtime="00:01:34.34" resultid="2380" heatid="4881" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="431" swimtime="00:01:06.49" resultid="2381" heatid="4932" lane="6" entrytime="00:01:08.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="400" swimtime="00:00:31.12" resultid="2382" heatid="5094" lane="6" entrytime="00:00:31.34" entrycourse="SCM" />
                <RESULT eventid="1301" points="262" swimtime="00:00:44.32" resultid="2383" heatid="5041" lane="3" entrytime="00:00:45.98" entrycourse="SCM" />
                <RESULT eventid="4411" points="320" swimtime="00:00:35.64" resultid="5392" heatid="4680" lane="6" />
                <RESULT eventid="5804" points="416" swimtime="00:00:30.71" resultid="10192" heatid="6054" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco" lastname="Vianna Almeida" birthdate="2014-12-16" gender="M" nation="BRA" license="410292" swrid="5740019" athleteid="3018" externalid="410292" level="CLBO">
              <RESULTS>
                <RESULT eventid="1089" points="71" swimtime="00:00:52.34" resultid="3019" heatid="4752" lane="1" />
                <RESULT eventid="1102" points="118" swimtime="00:00:44.97" resultid="3020" heatid="4815" lane="2" entrytime="00:00:50.21" entrycourse="SCM" />
                <RESULT eventid="1213" points="117" swimtime="00:01:52.72" resultid="3021" heatid="4948" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1249" points="97" swimtime="00:01:44.92" resultid="3022" heatid="4981" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1326" points="134" swimtime="00:00:48.66" resultid="3024" heatid="5131" lane="6" entrytime="00:00:52.62" entrycourse="SCM" />
                <RESULT eventid="4445" points="139" swimtime="00:00:48.10" resultid="10317" heatid="6034" lane="7" />
                <RESULT eventid="10329" points="129" swimtime="00:00:39.84" resultid="10462" heatid="10342" lane="3" entrytime="00:00:42.77" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT comment="SW 10.12 - Os pés perderam contato com a plataforma de partida antes que o colega de equipe anterior tocasse a borda." eventid="1115" status="DSQ" swimtime="00:04:41.86" resultid="3081" heatid="4871" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.91" />
                    <SPLIT distance="100" swimtime="00:01:14.77" />
                    <SPLIT distance="150" swimtime="00:01:48.16" />
                    <SPLIT distance="200" swimtime="00:02:24.28" />
                    <SPLIT distance="250" swimtime="00:02:55.59" />
                    <SPLIT distance="300" swimtime="00:03:33.26" />
                    <SPLIT distance="350" swimtime="00:04:16.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2767" number="1" />
                    <RELAYPOSITION athleteid="2594" number="2" />
                    <RELAYPOSITION athleteid="2524" number="3" />
                    <RELAYPOSITION athleteid="2426" number="4" />
                    <RELAYPOSITION athleteid="2309" number="5" />
                    <RELAYPOSITION athleteid="2356" number="6" />
                    <RELAYPOSITION athleteid="2183" number="7" />
                    <RELAYPOSITION athleteid="2211" number="8" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1339" points="247" swimtime="00:04:20.43" resultid="3082" heatid="5246" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.52" />
                    <SPLIT distance="100" swimtime="00:01:17.30" />
                    <SPLIT distance="150" swimtime="00:01:49.90" />
                    <SPLIT distance="200" swimtime="00:02:19.37" />
                    <SPLIT distance="250" swimtime="00:02:54.43" />
                    <SPLIT distance="300" swimtime="00:03:28.58" />
                    <SPLIT distance="350" swimtime="00:03:55.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2816" number="1" />
                    <RELAYPOSITION athleteid="2587" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2412" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="2344" number="4" reactiontime="0" />
                    <RELAYPOSITION athleteid="2475" number="5" reactiontime="0" />
                    <RELAYPOSITION athleteid="2489" number="6" reactiontime="0" />
                    <RELAYPOSITION athleteid="2183" number="7" reactiontime="0" />
                    <RELAYPOSITION athleteid="2608" number="8" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1115" points="252" swimtime="00:04:44.06" resultid="3085" heatid="4871" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.22" />
                    <SPLIT distance="100" swimtime="00:01:23.14" />
                    <SPLIT distance="150" swimtime="00:01:59.14" />
                    <SPLIT distance="200" swimtime="00:02:30.32" />
                    <SPLIT distance="250" swimtime="00:03:08.52" />
                    <SPLIT distance="300" swimtime="00:03:41.91" />
                    <SPLIT distance="350" swimtime="00:04:07.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3011" number="1" />
                    <RELAYPOSITION athleteid="2690" number="2" />
                    <RELAYPOSITION athleteid="2725" number="3" />
                    <RELAYPOSITION athleteid="3033" number="4" />
                    <RELAYPOSITION athleteid="2391" number="5" />
                    <RELAYPOSITION athleteid="2398" number="6" />
                    <RELAYPOSITION athleteid="2246" number="7" />
                    <RELAYPOSITION athleteid="2239" number="8" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1339" points="249" swimtime="00:04:19.86" resultid="3086" heatid="5246" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.52" />
                    <SPLIT distance="100" swimtime="00:01:15.42" />
                    <SPLIT distance="150" swimtime="00:01:45.77" />
                    <SPLIT distance="200" swimtime="00:02:16.71" />
                    <SPLIT distance="250" swimtime="00:02:53.25" />
                    <SPLIT distance="300" swimtime="00:03:25.75" />
                    <SPLIT distance="350" swimtime="00:03:52.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2928" number="1" />
                    <RELAYPOSITION athleteid="2690" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2552" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="2363" number="4" reactiontime="0" />
                    <RELAYPOSITION athleteid="2531" number="5" reactiontime="0" />
                    <RELAYPOSITION athleteid="2538" number="6" reactiontime="0" />
                    <RELAYPOSITION athleteid="2419" number="7" reactiontime="0" />
                    <RELAYPOSITION athleteid="2211" number="8" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;C&quot;" number="3">
              <RESULTS>
                <RESULT eventid="1115" points="232" status="EXH" swimtime="00:04:51.63" resultid="3089" heatid="4871" lane="6">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:01:48.37" />
                    <SPLIT distance="200" swimtime="00:02:24.13" />
                    <SPLIT distance="250" swimtime="00:02:59.36" />
                    <SPLIT distance="300" swimtime="00:03:43.49" />
                    <SPLIT distance="350" swimtime="00:04:23.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2746" number="1" />
                    <RELAYPOSITION athleteid="2412" number="2" />
                    <RELAYPOSITION athleteid="2316" number="3" />
                    <RELAYPOSITION athleteid="2879" number="4" />
                    <RELAYPOSITION athleteid="2337" number="5" />
                    <RELAYPOSITION athleteid="2517" number="6" />
                    <RELAYPOSITION athleteid="2288" number="7" />
                    <RELAYPOSITION athleteid="2232" number="8" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1339" points="215" status="EXH" swimtime="00:04:33.07" resultid="3090" heatid="5246" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                    <SPLIT distance="100" swimtime="00:01:16.35" />
                    <SPLIT distance="150" swimtime="00:01:48.00" />
                    <SPLIT distance="200" swimtime="00:02:19.38" />
                    <SPLIT distance="250" swimtime="00:03:01.18" />
                    <SPLIT distance="300" swimtime="00:03:36.54" />
                    <SPLIT distance="350" swimtime="00:04:04.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2886" number="1" />
                    <RELAYPOSITION athleteid="2594" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="2524" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="2725" number="4" reactiontime="0" />
                    <RELAYPOSITION athleteid="2503" number="5" reactiontime="0" />
                    <RELAYPOSITION athleteid="5256" number="6" reactiontime="0" />
                    <RELAYPOSITION athleteid="2246" number="7" reactiontime="0" />
                    <RELAYPOSITION athleteid="2288" number="8" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT comment="SW 10.12 - Os pés perderam contato com a plataforma de partida antes que o colega de equipe anterior tocasse a borda." eventid="1087" status="DSQ" swimtime="00:04:43.13" resultid="3079" heatid="4748" lane="5">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2823" number="1" />
                    <RELAYPOSITION athleteid="2566" number="2" />
                    <RELAYPOSITION athleteid="2963" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="2433" number="4" status="DSQ" />
                    <RELAYPOSITION athleteid="2377" number="5" status="DSQ" />
                    <RELAYPOSITION athleteid="2510" number="6" status="DSQ" />
                    <RELAYPOSITION athleteid="2302" number="7" status="DSQ" />
                    <RELAYPOSITION athleteid="2253" number="8" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1324" points="325" swimtime="00:04:28.92" resultid="3080" heatid="5123" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.70" />
                    <SPLIT distance="100" swimtime="00:01:15.66" />
                    <SPLIT distance="150" swimtime="00:01:47.06" />
                    <SPLIT distance="200" swimtime="00:02:19.85" />
                    <SPLIT distance="250" swimtime="00:02:54.19" />
                    <SPLIT distance="300" swimtime="00:03:29.36" />
                    <SPLIT distance="350" swimtime="00:03:58.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2809" number="1" />
                    <RELAYPOSITION athleteid="2566" number="2" />
                    <RELAYPOSITION athleteid="2704" number="3" />
                    <RELAYPOSITION athleteid="2454" number="4" />
                    <RELAYPOSITION athleteid="2496" number="5" />
                    <RELAYPOSITION athleteid="2615" number="6" />
                    <RELAYPOSITION athleteid="2190" number="7" />
                    <RELAYPOSITION athleteid="2281" number="8" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1087" points="333" swimtime="00:04:55.24" resultid="3083" heatid="4748" lane="4">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2788" number="1" />
                    <RELAYPOSITION athleteid="2844" number="2" />
                    <RELAYPOSITION athleteid="2858" number="3" />
                    <RELAYPOSITION athleteid="2461" number="4" />
                    <RELAYPOSITION athleteid="2330" number="5" />
                    <RELAYPOSITION athleteid="2323" number="6" />
                    <RELAYPOSITION athleteid="2281" number="7" />
                    <RELAYPOSITION athleteid="2601" number="8" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1324" points="294" swimtime="00:04:38.20" resultid="3084" heatid="5123" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.56" />
                    <SPLIT distance="100" swimtime="00:01:25.07" />
                    <SPLIT distance="150" swimtime="00:01:55.54" />
                    <SPLIT distance="200" swimtime="00:02:28.46" />
                    <SPLIT distance="250" swimtime="00:03:01.72" />
                    <SPLIT distance="300" swimtime="00:03:37.98" />
                    <SPLIT distance="350" swimtime="00:04:07.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2837" number="1" />
                    <RELAYPOSITION athleteid="2858" number="2" />
                    <RELAYPOSITION athleteid="2468" number="3" />
                    <RELAYPOSITION athleteid="2405" number="4" />
                    <RELAYPOSITION athleteid="2482" number="5" />
                    <RELAYPOSITION athleteid="2643" number="6" />
                    <RELAYPOSITION athleteid="2302" number="7" />
                    <RELAYPOSITION athleteid="2253" number="8" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;C&quot;" number="3">
              <RESULTS>
                <RESULT eventid="1087" points="328" status="EXH" swimtime="00:04:56.63" resultid="3087" heatid="4748" lane="2">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2760" number="1" />
                    <RELAYPOSITION athleteid="2669" number="2" />
                    <RELAYPOSITION athleteid="2440" number="3" />
                    <RELAYPOSITION athleteid="2545" number="4" />
                    <RELAYPOSITION athleteid="2370" number="5" />
                    <RELAYPOSITION athleteid="2384" number="6" />
                    <RELAYPOSITION athleteid="2190" number="7" />
                    <RELAYPOSITION athleteid="2197" number="8" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1324" points="273" status="EXH" swimtime="00:04:45.05" resultid="3088" heatid="5123" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="100" swimtime="00:01:06.22" />
                    <SPLIT distance="150" swimtime="00:01:37.08" />
                    <SPLIT distance="200" swimtime="00:02:13.99" />
                    <SPLIT distance="250" swimtime="00:02:48.35" />
                    <SPLIT distance="300" swimtime="00:03:19.52" />
                    <SPLIT distance="350" swimtime="00:03:47.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2774" number="1" />
                    <RELAYPOSITION athleteid="2718" number="2" />
                    <RELAYPOSITION athleteid="2384" number="3" />
                    <RELAYPOSITION athleteid="2942" number="4" />
                    <RELAYPOSITION athleteid="2711" number="5" />
                    <RELAYPOSITION athleteid="2963" number="6" />
                    <RELAYPOSITION athleteid="2197" number="7" />
                    <RELAYPOSITION athleteid="2447" number="8" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="3501" nation="BRA" region="PR" clubid="1924" swrid="93752" name="Ortega &amp; De Souza Jesus" shortname="Aquafoz">
          <ATHLETES>
            <ATHLETE firstname="Vitor" lastname="Gabriel Serighelli" birthdate="1999-03-12" gender="M" nation="BRA" license="121253" swrid="5596899" athleteid="1925" externalid="121253" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="578" swimtime="00:00:26.11" resultid="1926" heatid="4791" lane="4" entrytime="00:00:25.65" entrycourse="SCM" />
                <RESULT eventid="1105" points="460" swimtime="00:00:28.63" resultid="1927" heatid="4851" lane="4" entrytime="00:00:26.90" entrycourse="SCM" />
                <RESULT eventid="1249" points="504" swimtime="00:01:00.73" resultid="1928" heatid="4989" lane="3" entrytime="00:00:58.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="541" swimtime="00:00:24.73" resultid="1929" heatid="5226" lane="4" entrytime="00:00:24.36" entrycourse="SCM" />
                <RESULT eventid="1329" points="408" swimtime="00:00:33.63" resultid="1930" heatid="5156" lane="2" />
                <RESULT eventid="4423" points="546" swimtime="00:00:26.61" resultid="5722" heatid="4803" lane="2" />
                <RESULT eventid="4425" points="525" swimtime="00:00:26.95" resultid="5744" heatid="4809" lane="5" />
                <RESULT eventid="4429" points="481" swimtime="00:00:28.20" resultid="5772" heatid="4863" lane="2" />
                <RESULT eventid="4431" points="497" swimtime="00:00:27.91" resultid="5793" heatid="4869" lane="5" />
                <RESULT eventid="5807" points="392" swimtime="00:00:34.07" resultid="10153" heatid="6047" lane="6" />
                <RESULT eventid="5810" points="545" swimtime="00:00:24.68" resultid="10263" heatid="6031" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Victoria Portela" birthdate="2009-12-04" gender="F" nation="BRA" license="383047" swrid="5596945" athleteid="1951" externalid="383047" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="221" swimtime="00:00:40.27" resultid="1952" heatid="4673" lane="6" />
                <RESULT eventid="1077" points="210" swimtime="00:00:42.44" resultid="1953" heatid="4728" lane="2" entrytime="00:00:37.10" entrycourse="SCM" />
                <RESULT eventid="1143" points="372" swimtime="00:02:33.31" resultid="1954" heatid="4897" lane="2" entrytime="00:02:25.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.97" />
                    <SPLIT distance="100" swimtime="00:01:12.10" />
                    <SPLIT distance="150" swimtime="00:01:53.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="441" swimtime="00:01:05.98" resultid="1955" heatid="4939" lane="4" entrytime="00:01:05.03" entrycourse="SCM" />
                <RESULT eventid="1314" points="297" swimtime="00:00:34.35" resultid="1956" heatid="5103" lane="3" entrytime="00:00:29.33" entrycourse="SCM" />
                <RESULT eventid="1301" points="285" swimtime="00:00:43.10" resultid="1957" heatid="5051" lane="2" entrytime="00:00:40.42" entrycourse="SCM" />
                <RESULT eventid="4411" points="202" swimtime="00:00:41.55" resultid="5628" heatid="4687" lane="1" />
                <RESULT eventid="4413" points="283" swimtime="00:00:37.12" resultid="5645" heatid="4694" lane="4" />
                <RESULT eventid="4417" points="230" swimtime="00:00:41.20" resultid="5672" heatid="4738" lane="2" />
                <RESULT eventid="4419" points="302" swimtime="00:00:37.62" resultid="5690" heatid="4745" lane="5" />
                <RESULT eventid="5801" points="322" swimtime="00:00:41.37" resultid="10033" heatid="6075" lane="1" />
                <RESULT eventid="5804" points="422" swimtime="00:00:30.57" resultid="10072" heatid="6061" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruna" lastname="Mendes Portela" birthdate="2014-03-08" gender="F" nation="BRA" license="406656" swrid="5117156" athleteid="1997" externalid="406656" level="MRGA">
              <RESULTS>
                <RESULT eventid="1061" points="108" swimtime="00:00:51.11" resultid="1998" heatid="4652" lane="4" />
                <RESULT eventid="1074" points="133" swimtime="00:00:49.46" resultid="1999" heatid="4703" lane="3" />
                <RESULT eventid="1189" points="133" swimtime="00:01:38.38" resultid="2000" heatid="4936" lane="5" entrytime="00:01:50.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="125" swimtime="00:00:56.74" resultid="2001" heatid="5027" lane="5" entrytime="00:01:03.14" entrycourse="SCM" />
                <RESULT eventid="1311" points="155" swimtime="00:00:42.66" resultid="2002" heatid="5078" lane="3" entrytime="00:00:43.77" entrycourse="SCM" />
                <RESULT eventid="4433" points="125" swimtime="00:00:56.73" resultid="10010" heatid="6065" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Pires" birthdate="2011-04-09" gender="F" nation="BRA" license="383853" swrid="5596927" athleteid="1971" externalid="383853" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="197" swimtime="00:00:41.83" resultid="1972" heatid="4674" lane="5" />
                <RESULT eventid="1077" points="198" swimtime="00:00:43.32" resultid="1973" heatid="4724" lane="1" />
                <RESULT eventid="1129" points="215" swimtime="00:01:44.04" resultid="1974" heatid="4889" lane="3" entrytime="00:01:39.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="257" swimtime="00:00:36.02" resultid="1975" heatid="5099" lane="2" entrytime="00:00:36.93" entrycourse="SCM" />
                <RESULT eventid="1301" points="212" swimtime="00:00:47.53" resultid="1976" heatid="5050" lane="1" entrytime="00:00:47.87" entrycourse="SCM" />
                <RESULT eventid="4411" points="198" swimtime="00:00:41.77" resultid="5622" heatid="4683" lane="4" />
                <RESULT eventid="4413" points="179" swimtime="00:00:43.18" resultid="5641" heatid="4692" lane="6" />
                <RESULT eventid="4417" points="216" swimtime="00:00:42.06" resultid="5665" heatid="4734" lane="4" />
                <RESULT eventid="5801" points="220" swimtime="00:00:46.97" resultid="10025" heatid="6071" lane="3" />
                <RESULT eventid="5804" points="258" swimtime="00:00:36.01" resultid="10065" heatid="6057" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Marques Lima" birthdate="2010-04-30" gender="F" nation="BRA" license="383051" swrid="5596913" athleteid="1958" externalid="383051" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="367" swimtime="00:00:34.03" resultid="1959" heatid="4677" lane="5" entrytime="00:00:34.88" entrycourse="SCM" />
                <RESULT eventid="1077" points="293" swimtime="00:00:37.98" resultid="1960" heatid="4728" lane="4" entrytime="00:00:35.95" entrycourse="SCM" />
                <RESULT eventid="1119" points="334" swimtime="00:02:51.40" resultid="1961" heatid="4878" lane="4" entrytime="00:02:49.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.86" />
                    <SPLIT distance="100" swimtime="00:01:21.47" />
                    <SPLIT distance="150" swimtime="00:02:06.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1165" points="327" swimtime="00:01:19.65" resultid="1962" heatid="4917" lane="4" entrytime="00:01:18.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="343" swimtime="00:00:32.75" resultid="1963" heatid="5102" lane="5" entrytime="00:00:32.97" entrycourse="SCM" />
                <RESULT eventid="1301" points="211" swimtime="00:00:47.62" resultid="1964" heatid="5046" lane="3" />
                <RESULT eventid="4411" points="365" swimtime="00:00:34.10" resultid="5625" heatid="4685" lane="3" />
                <RESULT eventid="4413" points="340" swimtime="00:00:34.91" resultid="5644" heatid="4693" lane="6" />
                <RESULT eventid="4417" points="298" swimtime="00:00:37.77" resultid="5667" heatid="4736" lane="2" />
                <RESULT eventid="4419" points="328" swimtime="00:00:36.58" resultid="5687" heatid="4744" lane="5" />
                <RESULT eventid="5801" points="197" swimtime="00:00:48.68" resultid="10030" heatid="6073" lane="4" />
                <RESULT eventid="5804" points="338" swimtime="00:00:32.89" resultid="10068" heatid="6059" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Afonso Proteti" birthdate="2002-03-19" gender="M" nation="BRA" license="190464" swrid="5596865" athleteid="1938" externalid="190464" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="705" swimtime="00:00:24.43" resultid="1939" heatid="4791" lane="3" entrytime="00:00:24.70" entrycourse="SCM" />
                <RESULT eventid="1105" points="462" swimtime="00:00:28.58" resultid="1940" heatid="4851" lane="3" entrytime="00:00:26.75" entrycourse="SCM" />
                <RESULT comment="SW 8.5 - A cabeça não rompeu a superfície da água no ou antes do marco de 15m após o início ou a virada.  (Horário: 18:10), Na volta dos 25m." eventid="1237" status="DSQ" swimtime="00:00:54.66" resultid="1941" heatid="4977" lane="3" entrytime="00:00:55.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="555" swimtime="00:00:24.52" resultid="1942" heatid="5218" lane="4" />
                <RESULT eventid="1329" points="565" swimtime="00:00:30.17" resultid="1943" heatid="5160" lane="3" />
                <RESULT eventid="4423" points="590" swimtime="00:00:25.92" resultid="5721" heatid="4803" lane="1" />
                <RESULT eventid="4425" points="649" swimtime="00:00:25.12" resultid="5743" heatid="4809" lane="4" />
                <RESULT eventid="4429" points="491" swimtime="00:00:28.01" resultid="5771" heatid="4863" lane="1" />
                <RESULT eventid="4431" points="574" swimtime="00:00:26.60" resultid="5792" heatid="4869" lane="4" />
                <RESULT eventid="5807" points="560" swimtime="00:00:30.26" resultid="10148" heatid="6047" lane="1" />
                <RESULT eventid="5810" points="562" swimtime="00:00:24.42" resultid="10262" heatid="6031" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Mussi" birthdate="2006-12-31" gender="M" nation="BRA" license="370567" swrid="5596917" athleteid="1977" externalid="370567" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="443" swimtime="00:00:28.52" resultid="1978" heatid="4790" lane="3" entrytime="00:00:28.74" entrycourse="SCM" />
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="1979" heatid="4844" lane="5" />
                <RESULT eventid="1213" points="443" swimtime="00:01:12.49" resultid="1980" heatid="4959" lane="2" entrytime="00:01:10.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="393" swimtime="00:00:27.52" resultid="1981" heatid="5219" lane="6" />
                <RESULT eventid="1329" points="480" swimtime="00:00:31.86" resultid="1982" heatid="5165" lane="2" entrytime="00:00:31.45" entrycourse="SCM" />
                <RESULT eventid="4423" points="364" swimtime="00:00:30.45" resultid="5727" heatid="4803" lane="6" />
                <RESULT eventid="5807" points="487" swimtime="00:00:31.70" resultid="10150" heatid="6047" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luisa" lastname="Franco" birthdate="2010-06-09" gender="F" nation="BRA" license="383849" swrid="5596896" athleteid="1931" externalid="383849" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="435" swimtime="00:00:32.17" resultid="1932" heatid="4677" lane="4" entrytime="00:00:32.80" entrycourse="SCM" />
                <RESULT eventid="1077" points="312" swimtime="00:00:37.20" resultid="1933" heatid="4724" lane="3" />
                <RESULT eventid="1153" points="424" swimtime="00:01:11.93" resultid="1934" heatid="4903" lane="3" entrytime="00:01:15.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="380" swimtime="00:01:09.37" resultid="1935" heatid="4939" lane="1" entrytime="00:01:09.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="384" swimtime="00:00:31.54" resultid="1936" heatid="5102" lane="2" entrytime="00:00:32.32" entrycourse="SCM" />
                <RESULT eventid="1301" points="239" swimtime="00:00:45.71" resultid="1937" heatid="5048" lane="4" />
                <RESULT eventid="4411" points="384" swimtime="00:00:33.52" resultid="5623" heatid="4685" lane="1" />
                <RESULT eventid="4413" points="423" swimtime="00:00:32.46" resultid="5643" heatid="4693" lane="5" />
                <RESULT eventid="4417" points="229" swimtime="00:00:41.22" resultid="5666" heatid="4736" lane="1" />
                <RESULT eventid="5801" points="232" swimtime="00:00:46.17" resultid="10029" heatid="6073" lane="3" />
                <RESULT eventid="5804" points="370" swimtime="00:00:31.92" resultid="10067" heatid="6059" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kauan" lastname="Matheus Cunha" birthdate="2011-01-31" gender="M" nation="BRA" license="392834" swrid="5641770" athleteid="1983" externalid="392834" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="228" swimtime="00:00:35.60" resultid="1984" heatid="4788" lane="2" entrytime="00:00:36.83" entrycourse="SCM" />
                <RESULT eventid="1105" points="179" swimtime="00:00:39.17" resultid="1985" heatid="4848" lane="1" entrytime="00:00:45.04" entrycourse="SCM" />
                <RESULT eventid="1237" points="209" swimtime="00:01:20.48" resultid="1986" heatid="4976" lane="6" entrytime="00:01:46.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="274" swimtime="00:01:08.96" resultid="1987" heatid="5015" lane="3" entrytime="00:01:13.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="279" swimtime="00:00:30.83" resultid="1988" heatid="5222" lane="1" entrytime="00:00:32.42" entrycourse="SCM" />
                <RESULT eventid="1329" points="256" swimtime="00:00:39.27" resultid="1989" heatid="5161" lane="6" />
                <RESULT eventid="4423" points="221" swimtime="00:00:35.95" resultid="5712" heatid="4797" lane="6" />
                <RESULT eventid="5807" points="258" swimtime="00:00:39.19" resultid="10134" heatid="6041" lane="2" />
                <RESULT eventid="5810" points="288" swimtime="00:00:30.50" resultid="10250" heatid="6025" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Gustavo Cunha" birthdate="2011-01-31" gender="M" nation="BRA" license="392836" swrid="5641764" athleteid="1990" externalid="392836" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="175" swimtime="00:00:38.82" resultid="1991" heatid="4784" lane="4" />
                <RESULT eventid="1105" points="186" swimtime="00:00:38.73" resultid="1992" heatid="4842" lane="4" />
                <RESULT eventid="1227" points="267" swimtime="00:02:34.29" resultid="1993" heatid="5254" lane="1" entrytime="00:03:01.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                    <SPLIT distance="100" swimtime="00:01:14.23" />
                    <SPLIT distance="150" swimtime="00:01:54.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="274" swimtime="00:01:09.02" resultid="1994" heatid="5016" lane="2" entrytime="00:01:12.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="264" swimtime="00:00:31.42" resultid="1995" heatid="5222" lane="5" entrytime="00:00:32.08" entrycourse="SCM" />
                <RESULT eventid="1329" points="200" swimtime="00:00:42.65" resultid="1996" heatid="5163" lane="3" entrytime="00:00:43.60" entrycourse="SCM" />
                <RESULT eventid="5807" points="214" swimtime="00:00:41.67" resultid="10137" heatid="6041" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julio" lastname="Heck" birthdate="1998-02-15" gender="M" nation="BRA" license="185880" swrid="5596906" athleteid="1965" externalid="185880" level="MRGA">
              <RESULTS>
                <RESULT eventid="1092" points="451" swimtime="00:00:28.36" resultid="1966" heatid="4784" lane="6" />
                <RESULT eventid="1105" points="329" swimtime="00:00:32.00" resultid="1967" heatid="4851" lane="2" entrytime="00:00:29.95" entrycourse="SCM" />
                <RESULT eventid="1273" points="644" swimtime="00:00:51.91" resultid="1968" heatid="5018" lane="3" entrytime="00:00:51.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="618" swimtime="00:00:23.66" resultid="1969" heatid="5226" lane="3" entrytime="00:00:23.43" entrycourse="SCM" />
                <RESULT eventid="1329" points="276" swimtime="00:00:38.30" resultid="1970" heatid="5162" lane="6" />
                <RESULT eventid="4423" points="411" swimtime="00:00:29.24" resultid="5723" heatid="4803" lane="3" />
                <RESULT eventid="5810" points="591" swimtime="00:00:24.02" resultid="10261" heatid="6031" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Geórgia" lastname="Adeli Jesus" birthdate="2008-03-27" gender="F" nation="BRA" license="312649" swrid="5596864" athleteid="1944" externalid="312649" level="MRGA">
              <RESULTS>
                <RESULT eventid="1064" points="267" swimtime="00:00:37.84" resultid="1945" heatid="4673" lane="4" />
                <RESULT eventid="1077" points="244" swimtime="00:00:40.39" resultid="1946" heatid="4725" lane="1" />
                <RESULT eventid="1143" points="423" swimtime="00:02:26.94" resultid="1947" heatid="4897" lane="4" entrytime="00:02:24.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                    <SPLIT distance="100" swimtime="00:01:09.35" />
                    <SPLIT distance="150" swimtime="00:01:47.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1189" points="390" swimtime="00:01:08.76" resultid="1948" heatid="4939" lane="5" entrytime="00:01:08.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1314" points="293" swimtime="00:00:34.51" resultid="1949" heatid="5098" lane="1" />
                <RESULT eventid="1301" points="164" swimtime="00:00:51.75" resultid="1950" heatid="5046" lane="1" />
                <RESULT eventid="4411" points="230" swimtime="00:00:39.76" resultid="5631" heatid="4689" lane="2" />
                <RESULT eventid="4413" points="310" swimtime="00:00:36.01" resultid="5648" heatid="4695" lane="5" />
                <RESULT eventid="4417" points="255" swimtime="00:00:39.80" resultid="5674" heatid="4740" lane="2" />
                <RESULT eventid="4419" points="217" swimtime="00:00:42.00" resultid="5692" heatid="4746" lane="5" />
                <RESULT eventid="5801" points="157" swimtime="00:00:52.52" resultid="10038" heatid="6077" lane="3" />
                <RESULT eventid="5804" points="285" swimtime="00:00:34.83" resultid="10074" heatid="6063" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
